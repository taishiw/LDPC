/* */

module ctrl(/*AUTOARG*/
	    //Inputs
	    i_data,i_val,
	    //Outputs
	    estimate,o_val,clk,xrst,r_loop
	    );
   input [15:0] i_data;//雑音の付加されたデータ
   input 	     i_val;//入力のvalid信号
   output reg [399:0] estimate;//推定結果
   output 		   o_val;//出力のvalid信号
   input 		   clk;//クロック信号
   input 		   xrst;//リセット信号
   output reg [6:0] 	      r_loop;//繰り返し回数レジスタ
   //ステート情報
   parameter zStateInit=0;
   parameter zStateLambdaInit=1;
   parameter zStateBetaInit=2;
   parameter zStateRow=3;
   parameter zStateEstimate=4;
   parameter zStateColumn=5;
   
   reg [2:0] r_state;//ステートレジスタ
   
   reg [30:0] 			 r_counter;// カウンタ   
   reg [2:0] 			 i_init_row;//行処理の初期化信号
   reg [2:0] 			 i_init_column;//列処理の初期化信号
   
   wire 			 parity;//パリティビット
   
   wire [15:0]   w_i_data_row,w_i_data_column;//行処理，列処理それぞれの入力信号
   wire [15:0]   w_o_data_column,w_o_data_row;//行処理，列処理の出力信号
   reg 			   r_i_val_row,r_i_val_column;//行処理，列処理の入力のvalid信号
   wire 		   w_o_val_row,w_o_val_column;//行処理，列処理の出力のvalid信号
   wire 		   w_trans_row,w_trans_column,w_trans_lambdainit,w_trans_betainit,w_trans_estimate;//行処理，列処理の状態遷移
   wire signed [15:0] o_data_test_alpha,o_data_test_beta;
   wire signed [15:0] o_column_data;
   
   
   //sram関係
   
   //lambda
   wire 			   i_wen_lambda;
   wire [19:0] 			   i_waddr_lambda,i_raddr_lambda;
   wire [15:0] 	   i_wdata_lambda;
   wire [15:0] 	   o_rdata_lambda;

   //alpha
   wire 			   i_wen_alpha;
   wire [19:0] 			   i_waddr_alpha,i_raddr_alpha;
   wire [15:0] 	   i_wdata_alpha;
   wire [15:0] 	   o_rdata_alpha;

   //beta
   wire 			   i_wen_beta;
   wire [19:0] 			   i_waddr_beta,i_raddr_beta;
   wire [15:0] 	   i_wdata_beta;
   wire [15:0] 	   o_rdata_beta;
   
   
   assign w_trans_lambdainit = (r_state==zStateInit & i_val);

   assign w_trans_betainit = (r_state == zStateLambdaInit) & (r_counter == 399);
   //ステートが初期値のときvalid信号をうけたら，行処理にステートを移す
   assign w_trans_row = (r_state==zStateBetaInit & r_counter==800) | (r_state==zStateColumn & r_counter==1602);

   assign w_trans_estimate=  (r_state == zStateRow) & (r_counter == 2402) & w_o_val_row; 

   //ステートが行処理かつカウンタが行処理の最後の処理かつ行処理の出力valid信号が１のときステートを列処理に移す
   assign w_trans_column = (r_state == zStateEstimate) & (r_counter == 1201); 
   /*パリティビットを計算
    行を取り出し，検査行列を1が立っている列の推定結果の和を
    だして，すべての列の積をとる
    */ 
   assign parity=  /**/
		   (
		    /**/
		    estimate[274]^
	            /**/
		    estimate[198]^
	            /**/
		    estimate[197]^
	            /**/
       		    estimate[196] ==0) &
		   /**/
		   (
		    /**/
		    estimate[195]^
	            /**/
		    estimate[194]^
	            /**/
		    estimate[193]^
	            /**/
       		    estimate[192] ==0) &
		   /**/
		   (
		    /**/
		    estimate[191]^
	            /**/
		    estimate[190]^
	            /**/
		    estimate[189]^
	            /**/
       		    estimate[188] ==0) &
		   /**/
		   (
		    /**/
		    estimate[187]^
	            /**/
		    estimate[186]^
	            /**/
		    estimate[185]^
	            /**/
       		    estimate[184] ==0) &
		   /**/
		   (
		    /**/
		    estimate[183]^
	            /**/
		    estimate[182]^
	            /**/
		    estimate[181]^
	            /**/
       		    estimate[180] ==0) &
		   /**/
		   (
		    /**/
		    estimate[179]^
	            /**/
		    estimate[178]^
	            /**/
		    estimate[177]^
	            /**/
       		    estimate[176] ==0) &
		   /**/
		   (
		    /**/
		    estimate[175]^
	            /**/
		    estimate[174]^
	            /**/
		    estimate[173]^
	            /**/
       		    estimate[172] ==0) &
		   /**/
		   (
		    /**/
		    estimate[171]^
	            /**/
		    estimate[170]^
	            /**/
		    estimate[169]^
	            /**/
       		    estimate[168] ==0) &
		   /**/
		   (
		    /**/
		    estimate[167]^
	            /**/
		    estimate[166]^
	            /**/
		    estimate[165]^
	            /**/
       		    estimate[164] ==0) &
		   /**/
		   (
		    /**/
		    estimate[163]^
	            /**/
		    estimate[162]^
	            /**/
		    estimate[161]^
	            /**/
       		    estimate[160] ==0) &
		   /**/
		   (
		    /**/
		    estimate[159]^
	            /**/
		    estimate[158]^
	            /**/
		    estimate[157]^
	            /**/
       		    estimate[156] ==0) &
		   /**/
		   (
		    /**/
		    estimate[155]^
	            /**/
		    estimate[154]^
	            /**/
		    estimate[153]^
	            /**/
       		    estimate[152] ==0) &
		   /**/
		   (
		    /**/
		    estimate[390]^
	            /**/
		    estimate[151]^
	            /**/
		    estimate[150]^
	            /**/
       		    estimate[149] ==0) &
		   /**/
		   (
		    /**/
		    estimate[148]^
	            /**/
		    estimate[147]^
	            /**/
		    estimate[146]^
	            /**/
       		    estimate[145] ==0) &
		   /**/
		   (
		    /**/
		    estimate[144]^
	            /**/
		    estimate[143]^
	            /**/
		    estimate[142]^
	            /**/
       		    estimate[141] ==0) &
		   /**/
		   (
		    /**/
		    estimate[140]^
	            /**/
		    estimate[139]^
	            /**/
		    estimate[138]^
	            /**/
       		    estimate[137] ==0) &
		   /**/
		   (
		    /**/
		    estimate[338]^
	            /**/
		    estimate[136]^
	            /**/
		    estimate[135]^
	            /**/
       		    estimate[134] ==0) &
		   /**/
		   (
		    /**/
		    estimate[133]^
	            /**/
		    estimate[132]^
	            /**/
		    estimate[131]^
	            /**/
       		    estimate[130] ==0) &
		   /**/
		   (
		    /**/
		    estimate[370]^
	            /**/
		    estimate[129]^
	            /**/
		    estimate[128]^
	            /**/
       		    estimate[127] ==0) &
		   /**/
		   (
		    /**/
		    estimate[126]^
	            /**/
		    estimate[125]^
	            /**/
		    estimate[124]^
	            /**/
       		    estimate[123] ==0) &
		   /**/
		   (
		    /**/
		    estimate[122]^
	            /**/
		    estimate[121]^
	            /**/
		    estimate[120]^
	            /**/
       		    estimate[119] ==0) &
		   /**/
		   (
		    /**/
		    estimate[298]^
	            /**/
		    estimate[118]^
	            /**/
		    estimate[117]^
	            /**/
       		    estimate[116] ==0) &
		   /**/
		   (
		    /**/
		    estimate[386]^
	            /**/
		    estimate[115]^
	            /**/
		    estimate[114]^
	            /**/
       		    estimate[113] ==0) &
		   /**/
		   (
		    /**/
		    estimate[112]^
	            /**/
		    estimate[111]^
	            /**/
		    estimate[110]^
	            /**/
       		    estimate[109] ==0) &
		   /**/
		   (
		    /**/
		    estimate[346]^
	            /**/
		    estimate[345]^
	            /**/
		    estimate[108]^
	            /**/
       		    estimate[107] ==0) &
		   /**/
		   (
		    /**/
		    estimate[242]^
	            /**/
		    estimate[106]^
	            /**/
		    estimate[105]^
	            /**/
       		    estimate[104] ==0) &
		   /**/
		   (
		    /**/
		    estimate[103]^
	            /**/
		    estimate[102]^
	            /**/
		    estimate[101]^
	            /**/
       		    estimate[100] ==0) &
		   /**/
		   (
		    /**/
		    estimate[334]^
	            /**/
		    estimate[99]^
	            /**/
		    estimate[98]^
	            /**/
       		    estimate[97] ==0) &
		   /**/
		   (
		    /**/
		    estimate[394]^
	            /**/
		    estimate[226]^
	            /**/
		    estimate[96]^
	            /**/
       		    estimate[95] ==0) &
		   /**/
		   (
		    /**/
		    estimate[382]^
	            /**/
		    estimate[378]^
	            /**/
		    estimate[94]^
	            /**/
       		    estimate[93] ==0) &
		   /**/
		   (
		    /**/
		    estimate[366]^
	            /**/
		    estimate[358]^
	            /**/
		    estimate[350]^
	            /**/
       		    estimate[92] ==0) &
		   /**/
		   (
		    /**/
		    estimate[342]^
	            /**/
		    estimate[91]^
	            /**/
		    estimate[90]^
	            /**/
       		    estimate[89] ==0) &
		   /**/
		   (
		    /**/
		    estimate[330]^
	            /**/
		    estimate[314]^
	            /**/
		    estimate[302]^
	            /**/
       		    estimate[88] ==0) &
		   /**/
		   (
		    /**/
		    estimate[294]^
	            /**/
		    estimate[289]^
	            /**/
		    estimate[278]^
	            /**/
       		    estimate[87] ==0) &
		   /**/
		   (
		    /**/
		    estimate[270]^
	            /**/
		    estimate[266]^
	            /**/
		    estimate[258]^
	            /**/
       		    estimate[86] ==0) &
		   /**/
		   (
		    /**/
		    estimate[398]^
	            /**/
		    estimate[210]^
	            /**/
		    estimate[85]^
	            /**/
       		    estimate[84] ==0) &
		   /**/
		   (
		    /**/
		    estimate[383]^
	            /**/
		    estimate[83]^
	            /**/
		    estimate[82]^
	            /**/
       		    estimate[81] ==0) &
		   /**/
		   (
		    /**/
		    estimate[376]^
	            /**/
		    estimate[374]^
	            /**/
		    estimate[80]^
	            /**/
       		    estimate[79] ==0) &
		   /**/
		   (
		    /**/
		    estimate[369]^
	            /**/
		    estimate[362]^
	            /**/
		    estimate[78]^
	            /**/
       		    estimate[77] ==0) &
		   /**/
		   (
		    /**/
		    estimate[354]^
	            /**/
		    estimate[76]^
	            /**/
		    estimate[75]^
	            /**/
       		    estimate[74] ==0) &
		   /**/
		   (
		    /**/
		    estimate[73]^
	            /**/
		    estimate[72]^
	            /**/
		    estimate[71]^
	            /**/
       		    estimate[70] ==0) &
		   /**/
		   (
		    /**/
		    estimate[326]^
	            /**/
		    estimate[322]^
	            /**/
		    estimate[318]^
	            /**/
       		    estimate[69] ==0) &
		   /**/
		   (
		    /**/
		    estimate[310]^
	            /**/
		    estimate[308]^
	            /**/
		    estimate[306]^
	            /**/
       		    estimate[68] ==0) &
		   /**/
		   (
		    /**/
		    estimate[290]^
	            /**/
		    estimate[67]^
	            /**/
		    estimate[66]^
	            /**/
       		    estimate[65] ==0) &
		   /**/
		   (
		    /**/
		    estimate[286]^
	            /**/
		    estimate[282]^
	            /**/
		    estimate[64]^
	            /**/
       		    estimate[63] ==0) &
		   /**/
		   (
		    /**/
		    estimate[262]^
	            /**/
		    estimate[62]^
	            /**/
		    estimate[61]^
	            /**/
       		    estimate[60] ==0) &
		   /**/
		   (
		    /**/
		    estimate[254]^
	            /**/
		    estimate[250]^
	            /**/
		    estimate[246]^
	            /**/
       		    estimate[59] ==0) &
		   /**/
		   (
		    /**/
		    estimate[238]^
	            /**/
		    estimate[234]^
	            /**/
		    estimate[230]^
	            /**/
       		    estimate[58] ==0) &
		   /**/
		   (
		    /**/
		    estimate[222]^
	            /**/
		    estimate[218]^
	            /**/
		    estimate[214]^
	            /**/
       		    estimate[57] ==0) &
		   /**/
		   (
		    /**/
		    estimate[399]^
	            /**/
		    estimate[206]^
	            /**/
		    estimate[202]^
	            /**/
       		    estimate[56] ==0) &
		   /**/
		   (
		    /**/
		    estimate[397]^
	            /**/
		    estimate[396]^
	            /**/
		    estimate[395]^
	            /**/
       		    estimate[55] ==0) &
		   /**/
		   (
		    /**/
		    estimate[393]^
	            /**/
		    estimate[392]^
	            /**/
		    estimate[391]^
	            /**/
       		    estimate[54] ==0) &
		   /**/
		   (
		    /**/
		    estimate[389]^
	            /**/
		    estimate[388]^
	            /**/
		    estimate[387]^
	            /**/
       		    estimate[53] ==0) &
		   /**/
		   (
		    /**/
		    estimate[385]^
	            /**/
		    estimate[384]^
	            /**/
		    estimate[52]^
	            /**/
       		    estimate[51] ==0) &
		   /**/
		   (
		    /**/
		    estimate[381]^
	            /**/
		    estimate[380]^
	            /**/
		    estimate[379]^
	            /**/
       		    estimate[50] ==0) &
		   /**/
		   (
		    /**/
		    estimate[377]^
	            /**/
		    estimate[375]^
	            /**/
		    estimate[49]^
	            /**/
       		    estimate[48] ==0) &
		   /**/
		   (
		    /**/
		    estimate[373]^
	            /**/
		    estimate[372]^
	            /**/
		    estimate[371]^
	            /**/
       		    estimate[47] ==0) &
		   /**/
		   (
		    /**/
		    estimate[368]^
	            /**/
		    estimate[367]^
	            /**/
		    estimate[46]^
	            /**/
       		    estimate[45] ==0) &
		   /**/
		   (
		    /**/
		    estimate[365]^
	            /**/
		    estimate[364]^
	            /**/
		    estimate[363]^
	            /**/
       		    estimate[44] ==0) &
		   /**/
		   (
		    /**/
		    estimate[361]^
	            /**/
		    estimate[360]^
	            /**/
		    estimate[359]^
	            /**/
       		    estimate[43] ==0) &
		   /**/
		   (
		    /**/
		    estimate[357]^
	            /**/
		    estimate[356]^
	            /**/
		    estimate[355]^
	            /**/
       		    estimate[42] ==0) &
		   /**/
		   (
		    /**/
		    estimate[353]^
	            /**/
		    estimate[352]^
	            /**/
		    estimate[351]^
	            /**/
       		    estimate[41] ==0) &
		   /**/
		   (
		    /**/
		    estimate[349]^
	            /**/
		    estimate[348]^
	            /**/
		    estimate[347]^
	            /**/
       		    estimate[40] ==0) &
		   /**/
		   (
		    /**/
		    estimate[344]^
	            /**/
		    estimate[343]^
	            /**/
		    estimate[39]^
	            /**/
       		    estimate[38] ==0) &
		   /**/
		   (
		    /**/
		    estimate[341]^
	            /**/
		    estimate[340]^
	            /**/
		    estimate[339]^
	            /**/
       		    estimate[37] ==0) &
		   /**/
		   (
		    /**/
		    estimate[337]^
	            /**/
		    estimate[336]^
	            /**/
		    estimate[335]^
	            /**/
       		    estimate[36] ==0) &
		   /**/
		   (
		    /**/
		    estimate[333]^
	            /**/
		    estimate[332]^
	            /**/
		    estimate[331]^
	            /**/
       		    estimate[35] ==0) &
		   /**/
		   (
		    /**/
		    estimate[329]^
	            /**/
		    estimate[328]^
	            /**/
		    estimate[327]^
	            /**/
       		    estimate[34] ==0) &
		   /**/
		   (
		    /**/
		    estimate[325]^
	            /**/
		    estimate[324]^
	            /**/
		    estimate[323]^
	            /**/
       		    estimate[33] ==0) &
		   /**/
		   (
		    /**/
		    estimate[321]^
	            /**/
		    estimate[320]^
	            /**/
		    estimate[319]^
	            /**/
       		    estimate[32] ==0) &
		   /**/
		   (
		    /**/
		    estimate[317]^
	            /**/
		    estimate[316]^
	            /**/
		    estimate[315]^
	            /**/
       		    estimate[31] ==0) &
		   /**/
		   (
		    /**/
		    estimate[313]^
	            /**/
		    estimate[312]^
	            /**/
		    estimate[311]^
	            /**/
       		    estimate[30] ==0) &
		   /**/
		   (
		    /**/
		    estimate[309]^
	            /**/
		    estimate[307]^
	            /**/
		    estimate[29]^
	            /**/
       		    estimate[28] ==0) &
		   /**/
		   (
		    /**/
		    estimate[305]^
	            /**/
		    estimate[304]^
	            /**/
		    estimate[303]^
	            /**/
       		    estimate[27] ==0) &
		   /**/
		   (
		    /**/
		    estimate[301]^
	            /**/
		    estimate[300]^
	            /**/
		    estimate[299]^
	            /**/
       		    estimate[26] ==0) &
		   /**/
		   (
		    /**/
		    estimate[297]^
	            /**/
		    estimate[296]^
	            /**/
		    estimate[295]^
	            /**/
       		    estimate[25] ==0) &
		   /**/
		   (
		    /**/
		    estimate[293]^
	            /**/
		    estimate[292]^
	            /**/
		    estimate[291]^
	            /**/
       		    estimate[24] ==0) &
		   /**/
		   (
		    /**/
		    estimate[288]^
	            /**/
		    estimate[287]^
	            /**/
		    estimate[23]^
	            /**/
       		    estimate[22] ==0) &
		   /**/
		   (
		    /**/
		    estimate[285]^
	            /**/
		    estimate[284]^
	            /**/
		    estimate[283]^
	            /**/
       		    estimate[21] ==0) &
		   /**/
		   (
		    /**/
		    estimate[281]^
	            /**/
		    estimate[280]^
	            /**/
		    estimate[279]^
	            /**/
       		    estimate[20] ==0) &
		   /**/
		   (
		    /**/
		    estimate[277]^
	            /**/
		    estimate[276]^
	            /**/
		    estimate[275]^
	            /**/
       		    estimate[19] ==0) &
		   /**/
		   (
		    /**/
		    estimate[273]^
	            /**/
		    estimate[272]^
	            /**/
		    estimate[271]^
	            /**/
       		    estimate[18] ==0) &
		   /**/
		   (
		    /**/
		    estimate[269]^
	            /**/
		    estimate[268]^
	            /**/
		    estimate[267]^
	            /**/
       		    estimate[17] ==0) &
		   /**/
		   (
		    /**/
		    estimate[265]^
	            /**/
		    estimate[264]^
	            /**/
		    estimate[263]^
	            /**/
       		    estimate[16] ==0) &
		   /**/
		   (
		    /**/
		    estimate[261]^
	            /**/
		    estimate[260]^
	            /**/
		    estimate[259]^
	            /**/
       		    estimate[15] ==0) &
		   /**/
		   (
		    /**/
		    estimate[257]^
	            /**/
		    estimate[256]^
	            /**/
		    estimate[255]^
	            /**/
       		    estimate[14] ==0) &
		   /**/
		   (
		    /**/
		    estimate[253]^
	            /**/
		    estimate[252]^
	            /**/
		    estimate[251]^
	            /**/
       		    estimate[13] ==0) &
		   /**/
		   (
		    /**/
		    estimate[249]^
	            /**/
		    estimate[248]^
	            /**/
		    estimate[247]^
	            /**/
       		    estimate[12] ==0) &
		   /**/
		   (
		    /**/
		    estimate[245]^
	            /**/
		    estimate[244]^
	            /**/
		    estimate[243]^
	            /**/
       		    estimate[11] ==0) &
		   /**/
		   (
		    /**/
		    estimate[241]^
	            /**/
		    estimate[240]^
	            /**/
		    estimate[239]^
	            /**/
       		    estimate[10] ==0) &
		   /**/
		   (
		    /**/
		    estimate[237]^
	            /**/
		    estimate[236]^
	            /**/
		    estimate[235]^
	            /**/
       		    estimate[9] ==0) &
		   /**/
		   (
		    /**/
		    estimate[233]^
	            /**/
		    estimate[232]^
	            /**/
		    estimate[231]^
	            /**/
       		    estimate[8] ==0) &
		   /**/
		   (
		    /**/
		    estimate[229]^
	            /**/
		    estimate[228]^
	            /**/
		    estimate[227]^
	            /**/
       		    estimate[7] ==0) &
		   /**/
		   (
		    /**/
		    estimate[225]^
	            /**/
		    estimate[224]^
	            /**/
		    estimate[223]^
	            /**/
       		    estimate[6] ==0) &
		   /**/
		   (
		    /**/
		    estimate[221]^
	            /**/
		    estimate[220]^
	            /**/
		    estimate[219]^
	            /**/
       		    estimate[5] ==0) &
		   /**/
		   (
		    /**/
		    estimate[217]^
	            /**/
		    estimate[216]^
	            /**/
		    estimate[215]^
	            /**/
       		    estimate[4] ==0) &
		   /**/
		   (
		    /**/
		    estimate[213]^
	            /**/
		    estimate[212]^
	            /**/
		    estimate[211]^
	            /**/
       		    estimate[3] ==0) &
		   /**/
		   (
		    /**/
		    estimate[209]^
	            /**/
		    estimate[208]^
	            /**/
		    estimate[207]^
	            /**/
       		    estimate[2] ==0) &
		   /**/
		   (
		    /**/
		    estimate[205]^
	            /**/
		    estimate[204]^
	            /**/
		    estimate[203]^
	            /**/
       		    estimate[1] ==0) &
		   /**/
		   (
		    /**/
		    estimate[201]^
	            /**/
		    estimate[200]^
	            /**/
		    estimate[199]^
	            /**/
       		    estimate[0] ==0) &
		   /**/
		   (
		    /**/
		    estimate[325]^
	            /**/
		    estimate[264]^
	            /**/
		    estimate[221]^
	            /**/
       		    estimate[74] ==0) &
		   /**/
		   (
		    /**/
		    estimate[194]^
	            /**/
		    estimate[163]^
	            /**/
		    estimate[114]^
	            /**/
       		    estimate[64] ==0) &
		   /**/
		   (
		    /**/
		    estimate[377]^
	            /**/
		    estimate[317]^
	            /**/
		    estimate[65]^
	            /**/
       		    estimate[8] ==0) &
		   /**/
		   (
		    /**/
		    estimate[286]^
	            /**/
		    estimate[273]^
	            /**/
		    estimate[101]^
	            /**/
       		    estimate[70] ==0) &
		   /**/
		   (
		    /**/
		    estimate[391]^
	            /**/
		    estimate[330]^
	            /**/
		    estimate[104]^
	            /**/
       		    estimate[14] ==0) &
		   /**/
		   (
		    /**/
		    estimate[388]^
	            /**/
		    estimate[201]^
	            /**/
		    estimate[192]^
	            /**/
       		    estimate[67] ==0) &
		   /**/
		   (
		    /**/
		    estimate[210]^
	            /**/
		    estimate[141]^
	            /**/
		    estimate[128]^
	            /**/
       		    estimate[53] ==0) &
		   /**/
		   (
		    /**/
		    estimate[353]^
	            /**/
		    estimate[334]^
	            /**/
		    estimate[99]^
	            /**/
       		    estimate[52] ==0) &
		   /**/
		   (
		    /**/
		    estimate[347]^
	            /**/
		    estimate[298]^
	            /**/
		    estimate[189]^
	            /**/
       		    estimate[23] ==0) &
		   /**/
		   (
		    /**/
		    estimate[362]^
	            /**/
		    estimate[289]^
	            /**/
		    estimate[203]^
	            /**/
       		    estimate[142] ==0) &
		   /**/
		   (
		    /**/
		    estimate[238]^
	            /**/
		    estimate[122]^
	            /**/
		    estimate[87]^
	            /**/
       		    estimate[43] ==0) &
		   /**/
		   (
		    /**/
		    estimate[301]^
	            /**/
		    estimate[287]^
	            /**/
		    estimate[225]^
	            /**/
       		    estimate[82] ==0) &
		   /**/
		   (
		    /**/
		    estimate[338]^
	            /**/
		    estimate[311]^
	            /**/
		    estimate[269]^
	            /**/
       		    estimate[149] ==0) &
		   /**/
		   (
		    /**/
		    estimate[268]^
	            /**/
		    estimate[200]^
	            /**/
		    estimate[22]^
	            /**/
       		    estimate[0] ==0) &
		   /**/
		   (
		    /**/
		    estimate[335]^
	            /**/
		    estimate[297]^
	            /**/
		    estimate[75]^
	            /**/
       		    estimate[31] ==0) &
		   /**/
		   (
		    /**/
		    estimate[145]^
	            /**/
		    estimate[56]^
	            /**/
		    estimate[40]^
	            /**/
       		    estimate[27] ==0) &
		   /**/
		   (
		    /**/
		    estimate[389]^
	            /**/
		    estimate[369]^
	            /**/
		    estimate[219]^
	            /**/
       		    estimate[156] ==0) &
		   /**/
		   (
		    /**/
		    estimate[294]^
	            /**/
		    estimate[171]^
	            /**/
		    estimate[68]^
	            /**/
       		    estimate[34] ==0) &
		   /**/
		   (
		    /**/
		    estimate[381]^
	            /**/
		    estimate[320]^
	            /**/
		    estimate[173]^
	            /**/
       		    estimate[103] ==0) &
		   /**/
		   (
		    /**/
		    estimate[386]^
	            /**/
		    estimate[249]^
	            /**/
		    estimate[205]^
	            /**/
       		    estimate[119] ==0) &
		   /**/
		   (
		    /**/
		    estimate[303]^
	            /**/
		    estimate[263]^
	            /**/
		    estimate[204]^
	            /**/
       		    estimate[84] ==0) &
		   /**/
		   (
		    /**/
		    estimate[280]^
	            /**/
		    estimate[270]^
	            /**/
		    estimate[147]^
	            /**/
       		    estimate[46] ==0) &
		   /**/
		   (
		    /**/
		    estimate[226]^
	            /**/
		    estimate[197]^
	            /**/
		    estimate[176]^
	            /**/
       		    estimate[10] ==0) &
		   /**/
		   (
		    /**/
		    estimate[349]^
	            /**/
		    estimate[262]^
	            /**/
		    estimate[170]^
	            /**/
       		    estimate[127] ==0) &
		   /**/
		   (
		    /**/
		    estimate[383]^
	            /**/
		    estimate[359]^
	            /**/
		    estimate[313]^
	            /**/
       		    estimate[106] ==0) &
		   /**/
		   (
		    /**/
		    estimate[300]^
	            /**/
		    estimate[178]^
	            /**/
		    estimate[155]^
	            /**/
       		    estimate[132] ==0) &
		   /**/
		   (
		    /**/
		    estimate[361]^
	            /**/
		    estimate[304]^
	            /**/
		    estimate[215]^
	            /**/
       		    estimate[72] ==0) &
		   /**/
		   (
		    /**/
		    estimate[346]^
	            /**/
		    estimate[193]^
	            /**/
		    estimate[157]^
	            /**/
       		    estimate[151] ==0) &
		   /**/
		   (
		    /**/
		    estimate[396]^
	            /**/
		    estimate[327]^
	            /**/
		    estimate[161]^
	            /**/
       		    estimate[16] ==0) &
		   /**/
		   (
		    /**/
		    estimate[354]^
	            /**/
		    estimate[187]^
	            /**/
		    estimate[148]^
	            /**/
       		    estimate[20] ==0) &
		   /**/
		   (
		    /**/
		    estimate[231]^
	            /**/
		    estimate[217]^
	            /**/
		    estimate[100]^
	            /**/
       		    estimate[7] ==0) &
		   /**/
		   (
		    /**/
		    estimate[321]^
	            /**/
		    estimate[209]^
	            /**/
		    estimate[113]^
	            /**/
       		    estimate[15] ==0) &
		   /**/
		   (
		    /**/
		    estimate[340]^
	            /**/
		    estimate[332]^
	            /**/
		    estimate[212]^
	            /**/
       		    estimate[45] ==0) &
		   /**/
		   (
		    /**/
		    estimate[310]^
	            /**/
		    estimate[291]^
	            /**/
		    estimate[125]^
	            /**/
       		    estimate[24] ==0) &
		   /**/
		   (
		    /**/
		    estimate[246]^
	            /**/
		    estimate[186]^
	            /**/
		    estimate[153]^
	            /**/
       		    estimate[1] ==0) &
		   /**/
		   (
		    /**/
		    estimate[363]^
	            /**/
		    estimate[138]^
	            /**/
		    estimate[129]^
	            /**/
       		    estimate[116] ==0) &
		   /**/
		   (
		    /**/
		    estimate[281]^
	            /**/
		    estimate[255]^
	            /**/
		    estimate[248]^
	            /**/
       		    estimate[28] ==0) &
		   /**/
		   (
		    /**/
		    estimate[323]^
	            /**/
		    estimate[292]^
	            /**/
		    estimate[107]^
	            /**/
       		    estimate[69] ==0) &
		   /**/
		   (
		    /**/
		    estimate[374]^
	            /**/
		    estimate[364]^
	            /**/
		    estimate[185]^
	            /**/
       		    estimate[105] ==0) &
		   /**/
		   (
		    /**/
		    estimate[350]^
	            /**/
		    estimate[237]^
	            /**/
		    estimate[175]^
	            /**/
       		    estimate[17] ==0) &
		   /**/
		   (
		    /**/
		    estimate[394]^
	            /**/
		    estimate[190]^
	            /**/
		    estimate[126]^
	            /**/
       		    estimate[55] ==0) &
		   /**/
		   (
		    /**/
		    estimate[365]^
	            /**/
		    estimate[274]^
	            /**/
		    estimate[198]^
	            /**/
       		    estimate[80] ==0) &
		   /**/
		   (
		    /**/
		    estimate[259]^
	            /**/
		    estimate[253]^
	            /**/
		    estimate[79]^
	            /**/
       		    estimate[11] ==0) &
		   /**/
		   (
		    /**/
		    estimate[380]^
	            /**/
		    estimate[216]^
	            /**/
		    estimate[89]^
	            /**/
       		    estimate[26] ==0) &
		   /**/
		   (
		    /**/
		    estimate[351]^
	            /**/
		    estimate[342]^
	            /**/
		    estimate[229]^
	            /**/
       		    estimate[165] ==0) &
		   /**/
		   (
		    /**/
		    estimate[283]^
	            /**/
		    estimate[160]^
	            /**/
		    estimate[49]^
	            /**/
       		    estimate[35] ==0) &
		   /**/
		   (
		    /**/
		    estimate[367]^
	            /**/
		    estimate[272]^
	            /**/
		    estimate[247]^
	            /**/
       		    estimate[71] ==0) &
		   /**/
		   (
		    /**/
		    estimate[257]^
	            /**/
		    estimate[211]^
	            /**/
		    estimate[39]^
	            /**/
       		    estimate[3] ==0) &
		   /**/
		   (
		    /**/
		    estimate[241]^
	            /**/
		    estimate[181]^
	            /**/
		    estimate[133]^
	            /**/
       		    estimate[47] ==0) &
		   /**/
		   (
		    /**/
		    estimate[233]^
	            /**/
		    estimate[150]^
	            /**/
		    estimate[123]^
	            /**/
       		    estimate[76] ==0) &
		   /**/
		   (
		    /**/
		    estimate[356]^
	            /**/
		    estimate[202]^
	            /**/
		    estimate[180]^
	            /**/
       		    estimate[109] ==0) &
		   /**/
		   (
		    /**/
		    estimate[385]^
	            /**/
		    estimate[168]^
	            /**/
		    estimate[121]^
	            /**/
       		    estimate[12] ==0) &
		   /**/
		   (
		    /**/
		    estimate[337]^
	            /**/
		    estimate[277]^
	            /**/
		    estimate[256]^
	            /**/
       		    estimate[158] ==0) &
		   /**/
		   (
		    /**/
		    estimate[319]^
	            /**/
		    estimate[245]^
	            /**/
		    estimate[73]^
	            /**/
       		    estimate[5] ==0) &
		   /**/
		   (
		    /**/
		    estimate[232]^
	            /**/
		    estimate[228]^
	            /**/
		    estimate[207]^
	            /**/
       		    estimate[124] ==0) &
		   /**/
		   (
		    /**/
		    estimate[392]^
	            /**/
		    estimate[307]^
	            /**/
		    estimate[243]^
	            /**/
       		    estimate[60] ==0) &
		   /**/
		   (
		    /**/
		    estimate[384]^
	            /**/
		    estimate[329]^
	            /**/
		    estimate[98]^
	            /**/
       		    estimate[85] ==0) &
		   /**/
		   (
		    /**/
		    estimate[279]^
	            /**/
		    estimate[254]^
	            /**/
		    estimate[239]^
	            /**/
       		    estimate[62] ==0) &
		   /**/
		   (
		    /**/
		    estimate[348]^
	            /**/
		    estimate[267]^
	            /**/
		    estimate[261]^
	            /**/
       		    estimate[172] ==0) &
		   /**/
		   (
		    /**/
		    estimate[395]^
	            /**/
		    estimate[235]^
	            /**/
		    estimate[139]^
	            /**/
       		    estimate[108] ==0) &
		   /**/
		   (
		    /**/
		    estimate[315]^
	            /**/
		    estimate[227]^
	            /**/
		    estimate[191]^
	            /**/
       		    estimate[166] ==0) &
		   /**/
		   (
		    /**/
		    estimate[378]^
	            /**/
		    estimate[276]^
	            /**/
		    estimate[182]^
	            /**/
       		    estimate[96] ==0) &
		   /**/
		   (
		    /**/
		    estimate[293]^
	            /**/
		    estimate[102]^
	            /**/
		    estimate[58]^
	            /**/
       		    estimate[2] ==0) &
		   /**/
		   (
		    /**/
		    estimate[244]^
	            /**/
		    estimate[199]^
	            /**/
		    estimate[111]^
	            /**/
       		    estimate[36] ==0) &
		   /**/
		   (
		    /**/
		    estimate[370]^
	            /**/
		    estimate[188]^
	            /**/
		    estimate[137]^
	            /**/
       		    estimate[21] ==0) &
		   /**/
		   (
		    /**/
		    estimate[345]^
	            /**/
		    estimate[271]^
	            /**/
		    estimate[266]^
	            /**/
       		    estimate[130] ==0) &
		   /**/
		   (
		    /**/
		    estimate[393]^
	            /**/
		    estimate[331]^
	            /**/
		    estimate[179]^
	            /**/
       		    estimate[37] ==0) &
		   /**/
		   (
		    /**/
		    estimate[360]^
	            /**/
		    estimate[120]^
	            /**/
		    estimate[41]^
	            /**/
       		    estimate[32] ==0) &
		   /**/
		   (
		    /**/
		    estimate[344]^
	            /**/
		    estimate[295]^
	            /**/
		    estimate[284]^
	            /**/
       		    estimate[136] ==0) &
		   /**/
		   (
		    /**/
		    estimate[375]^
	            /**/
		    estimate[234]^
	            /**/
		    estimate[196]^
	            /**/
       		    estimate[97] ==0) &
		   /**/
		   (
		    /**/
		    estimate[305]^
	            /**/
		    estimate[51]^
	            /**/
		    estimate[6]^
	            /**/
       		    estimate[4] ==0) &
		   /**/
		   (
		    /**/
		    estimate[282]^
	            /**/
		    estimate[224]^
	            /**/
		    estimate[77]^
	            /**/
       		    estimate[18] ==0) &
		   /**/
		   (
		    /**/
		    estimate[372]^
	            /**/
		    estimate[368]^
	            /**/
		    estimate[144]^
	            /**/
       		    estimate[33] ==0) &
		   /**/
		   (
		    /**/
		    estimate[275]^
	            /**/
		    estimate[236]^
	            /**/
		    estimate[131]^
	            /**/
       		    estimate[9] ==0) &
		   /**/
		   (
		    /**/
		    estimate[357]^
	            /**/
		    estimate[220]^
	            /**/
		    estimate[112]^
	            /**/
       		    estimate[78] ==0) &
		   /**/
		   (
		    /**/
		    estimate[328]^
	            /**/
		    estimate[290]^
	            /**/
		    estimate[242]^
	            /**/
       		    estimate[115] ==0) &
		   /**/
		   (
		    /**/
		    estimate[371]^
	            /**/
		    estimate[230]^
	            /**/
		    estimate[174]^
	            /**/
       		    estimate[167] ==0) &
		   /**/
		   (
		    /**/
		    estimate[318]^
	            /**/
		    estimate[250]^
	            /**/
		    estimate[110]^
	            /**/
       		    estimate[25] ==0) &
		   /**/
		   (
		    /**/
		    estimate[358]^
	            /**/
		    estimate[278]^
	            /**/
		    estimate[169]^
	            /**/
       		    estimate[94] ==0) &
		   /**/
		   (
		    /**/
		    estimate[366]^
	            /**/
		    estimate[308]^
	            /**/
		    estimate[285]^
	            /**/
       		    estimate[183] ==0) &
		   /**/
		   (
		    /**/
		    estimate[265]^
	            /**/
		    estimate[260]^
	            /**/
		    estimate[66]^
	            /**/
       		    estimate[42] ==0) &
		   /**/
		   (
		    /**/
		    estimate[373]^
	            /**/
		    estimate[352]^
	            /**/
		    estimate[222]^
	            /**/
       		    estimate[140] ==0) &
		   /**/
		   (
		    /**/
		    estimate[339]^
	            /**/
		    estimate[296]^
	            /**/
		    estimate[81]^
	            /**/
       		    estimate[61] ==0) &
		   /**/
		   (
		    /**/
		    estimate[397]^
	            /**/
		    estimate[258]^
	            /**/
		    estimate[146]^
	            /**/
       		    estimate[117] ==0) &
		   /**/
		   (
		    /**/
		    estimate[306]^
	            /**/
		    estimate[177]^
	            /**/
		    estimate[86]^
	            /**/
       		    estimate[83] ==0) &
		   /**/
		   (
		    /**/
		    estimate[382]^
	            /**/
		    estimate[223]^
	            /**/
		    estimate[154]^
	            /**/
       		    estimate[29] ==0) &
		   /**/
		   (
		    /**/
		    estimate[312]^
	            /**/
		    estimate[299]^
	            /**/
		    estimate[159]^
	            /**/
       		    estimate[134] ==0) &
		   /**/
		   (
		    /**/
		    estimate[336]^
	            /**/
		    estimate[322]^
	            /**/
		    estimate[118]^
	            /**/
       		    estimate[50] ==0) &
		   /**/
		   (
		    /**/
		    estimate[341]^
	            /**/
		    estimate[333]^
	            /**/
		    estimate[251]^
	            /**/
       		    estimate[93] ==0) &
		   /**/
		   (
		    /**/
		    estimate[302]^
	            /**/
		    estimate[91]^
	            /**/
		    estimate[57]^
	            /**/
       		    estimate[44] ==0) &
		   /**/
		   (
		    /**/
		    estimate[240]^
	            /**/
		    estimate[208]^
	            /**/
		    estimate[63]^
	            /**/
       		    estimate[54] ==0) &
		   /**/
		   (
		    /**/
		    estimate[355]^
	            /**/
		    estimate[326]^
	            /**/
		    estimate[184]^
	            /**/
       		    estimate[90] ==0) &
		   /**/
		   (
		    /**/
		    estimate[343]^
	            /**/
		    estimate[324]^
	            /**/
		    estimate[164]^
	            /**/
       		    estimate[92] ==0) &
		   /**/
		   (
		    /**/
		    estimate[398]^
	            /**/
		    estimate[376]^
	            /**/
		    estimate[135]^
	            /**/
       		    estimate[13] ==0) &
		   /**/
		   (
		    /**/
		    estimate[379]^
	            /**/
		    estimate[309]^
	            /**/
		    estimate[252]^
	            /**/
       		    estimate[162] ==0) &
		   /**/
		   (
		    /**/
		    estimate[288]^
	            /**/
		    estimate[213]^
	            /**/
		    estimate[48]^
	            /**/
       		    estimate[30] ==0) &
		   /**/
		   (
		    /**/
		    estimate[399]^
	            /**/
		    estimate[214]^
	            /**/
		    estimate[152]^
	            /**/
       		    estimate[59] ==0) &
		   /**/
		   (
		    /**/
		    estimate[387]^
	            /**/
		    estimate[95]^
	            /**/
		    estimate[38]^
	            /**/
       		    estimate[19] ==0) &
		   /**/
		   (
		    /**/
		    estimate[390]^
	            /**/
		    estimate[206]^
	            /**/
		    estimate[195]^
	            /**/
       		    estimate[88] ==0) &
		   /**/
		   (
		    /**/
		    estimate[316]^
		    /**/
		    estimate[314]^
		    /**/
		    estimate[218]^
		    /**/
		    estimate[143] ==0);
   
   /*    推定結果を計算
    列を取り出し，検査行列で1が立っている行のαとその列のλの和をとり，
    0より大きければ0，小さければ1とする
    */
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[399] <= 0;
	else if(r_state == zStateEstimate & r_counter == 4)
	  estimate[399] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[399] <=  estimate[399];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[398] <= 0;
	else if(r_state == zStateEstimate & r_counter == 7)
	  estimate[398] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[398] <=  estimate[398];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[397] <= 0;
	else if(r_state == zStateEstimate & r_counter == 10)
	  estimate[397] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[397] <=  estimate[397];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[396] <= 0;
	else if(r_state == zStateEstimate & r_counter == 13)
	  estimate[396] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[396] <=  estimate[396];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[395] <= 0;
	else if(r_state == zStateEstimate & r_counter == 16)
	  estimate[395] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[395] <=  estimate[395];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[394] <= 0;
	else if(r_state == zStateEstimate & r_counter == 19)
	  estimate[394] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[394] <=  estimate[394];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[393] <= 0;
	else if(r_state == zStateEstimate & r_counter == 22)
	  estimate[393] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[393] <=  estimate[393];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[392] <= 0;
	else if(r_state == zStateEstimate & r_counter == 25)
	  estimate[392] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[392] <=  estimate[392];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[391] <= 0;
	else if(r_state == zStateEstimate & r_counter == 28)
	  estimate[391] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[391] <=  estimate[391];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[390] <= 0;
	else if(r_state == zStateEstimate & r_counter == 31)
	  estimate[390] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[390] <=  estimate[390];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[389] <= 0;
	else if(r_state == zStateEstimate & r_counter == 34)
	  estimate[389] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[389] <=  estimate[389];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[388] <= 0;
	else if(r_state == zStateEstimate & r_counter == 37)
	  estimate[388] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[388] <=  estimate[388];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[387] <= 0;
	else if(r_state == zStateEstimate & r_counter == 40)
	  estimate[387] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[387] <=  estimate[387];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[386] <= 0;
	else if(r_state == zStateEstimate & r_counter == 43)
	  estimate[386] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[386] <=  estimate[386];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[385] <= 0;
	else if(r_state == zStateEstimate & r_counter == 46)
	  estimate[385] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[385] <=  estimate[385];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[384] <= 0;
	else if(r_state == zStateEstimate & r_counter == 49)
	  estimate[384] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[384] <=  estimate[384];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[383] <= 0;
	else if(r_state == zStateEstimate & r_counter == 52)
	  estimate[383] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[383] <=  estimate[383];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[382] <= 0;
	else if(r_state == zStateEstimate & r_counter == 55)
	  estimate[382] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[382] <=  estimate[382];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[381] <= 0;
	else if(r_state == zStateEstimate & r_counter == 58)
	  estimate[381] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[381] <=  estimate[381];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[380] <= 0;
	else if(r_state == zStateEstimate & r_counter == 61)
	  estimate[380] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[380] <=  estimate[380];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[379] <= 0;
	else if(r_state == zStateEstimate & r_counter == 64)
	  estimate[379] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[379] <=  estimate[379];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[378] <= 0;
	else if(r_state == zStateEstimate & r_counter == 67)
	  estimate[378] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[378] <=  estimate[378];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[377] <= 0;
	else if(r_state == zStateEstimate & r_counter == 70)
	  estimate[377] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[377] <=  estimate[377];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[376] <= 0;
	else if(r_state == zStateEstimate & r_counter == 73)
	  estimate[376] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[376] <=  estimate[376];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[375] <= 0;
	else if(r_state == zStateEstimate & r_counter == 76)
	  estimate[375] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[375] <=  estimate[375];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[374] <= 0;
	else if(r_state == zStateEstimate & r_counter == 79)
	  estimate[374] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[374] <=  estimate[374];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[373] <= 0;
	else if(r_state == zStateEstimate & r_counter == 82)
	  estimate[373] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[373] <=  estimate[373];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[372] <= 0;
	else if(r_state == zStateEstimate & r_counter == 85)
	  estimate[372] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[372] <=  estimate[372];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[371] <= 0;
	else if(r_state == zStateEstimate & r_counter == 88)
	  estimate[371] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[371] <=  estimate[371];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[370] <= 0;
	else if(r_state == zStateEstimate & r_counter == 91)
	  estimate[370] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[370] <=  estimate[370];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[369] <= 0;
	else if(r_state == zStateEstimate & r_counter == 94)
	  estimate[369] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[369] <=  estimate[369];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[368] <= 0;
	else if(r_state == zStateEstimate & r_counter == 97)
	  estimate[368] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[368] <=  estimate[368];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[367] <= 0;
	else if(r_state == zStateEstimate & r_counter == 100)
	  estimate[367] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[367] <=  estimate[367];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[366] <= 0;
	else if(r_state == zStateEstimate & r_counter == 103)
	  estimate[366] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[366] <=  estimate[366];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[365] <= 0;
	else if(r_state == zStateEstimate & r_counter == 106)
	  estimate[365] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[365] <=  estimate[365];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[364] <= 0;
	else if(r_state == zStateEstimate & r_counter == 109)
	  estimate[364] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[364] <=  estimate[364];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[363] <= 0;
	else if(r_state == zStateEstimate & r_counter == 112)
	  estimate[363] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[363] <=  estimate[363];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[362] <= 0;
	else if(r_state == zStateEstimate & r_counter == 115)
	  estimate[362] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[362] <=  estimate[362];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[361] <= 0;
	else if(r_state == zStateEstimate & r_counter == 118)
	  estimate[361] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[361] <=  estimate[361];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[360] <= 0;
	else if(r_state == zStateEstimate & r_counter == 121)
	  estimate[360] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[360] <=  estimate[360];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[359] <= 0;
	else if(r_state == zStateEstimate & r_counter == 124)
	  estimate[359] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[359] <=  estimate[359];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[358] <= 0;
	else if(r_state == zStateEstimate & r_counter == 127)
	  estimate[358] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[358] <=  estimate[358];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[357] <= 0;
	else if(r_state == zStateEstimate & r_counter == 130)
	  estimate[357] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[357] <=  estimate[357];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[356] <= 0;
	else if(r_state == zStateEstimate & r_counter == 133)
	  estimate[356] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[356] <=  estimate[356];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[355] <= 0;
	else if(r_state == zStateEstimate & r_counter == 136)
	  estimate[355] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[355] <=  estimate[355];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[354] <= 0;
	else if(r_state == zStateEstimate & r_counter == 139)
	  estimate[354] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[354] <=  estimate[354];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[353] <= 0;
	else if(r_state == zStateEstimate & r_counter == 142)
	  estimate[353] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[353] <=  estimate[353];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[352] <= 0;
	else if(r_state == zStateEstimate & r_counter == 145)
	  estimate[352] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[352] <=  estimate[352];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[351] <= 0;
	else if(r_state == zStateEstimate & r_counter == 148)
	  estimate[351] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[351] <=  estimate[351];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[350] <= 0;
	else if(r_state == zStateEstimate & r_counter == 151)
	  estimate[350] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[350] <=  estimate[350];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[349] <= 0;
	else if(r_state == zStateEstimate & r_counter == 154)
	  estimate[349] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[349] <=  estimate[349];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[348] <= 0;
	else if(r_state == zStateEstimate & r_counter == 157)
	  estimate[348] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[348] <=  estimate[348];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[347] <= 0;
	else if(r_state == zStateEstimate & r_counter == 160)
	  estimate[347] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[347] <=  estimate[347];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[346] <= 0;
	else if(r_state == zStateEstimate & r_counter == 163)
	  estimate[346] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[346] <=  estimate[346];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[345] <= 0;
	else if(r_state == zStateEstimate & r_counter == 166)
	  estimate[345] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[345] <=  estimate[345];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[344] <= 0;
	else if(r_state == zStateEstimate & r_counter == 169)
	  estimate[344] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[344] <=  estimate[344];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[343] <= 0;
	else if(r_state == zStateEstimate & r_counter == 172)
	  estimate[343] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[343] <=  estimate[343];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[342] <= 0;
	else if(r_state == zStateEstimate & r_counter == 175)
	  estimate[342] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[342] <=  estimate[342];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[341] <= 0;
	else if(r_state == zStateEstimate & r_counter == 178)
	  estimate[341] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[341] <=  estimate[341];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[340] <= 0;
	else if(r_state == zStateEstimate & r_counter == 181)
	  estimate[340] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[340] <=  estimate[340];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[339] <= 0;
	else if(r_state == zStateEstimate & r_counter == 184)
	  estimate[339] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[339] <=  estimate[339];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[338] <= 0;
	else if(r_state == zStateEstimate & r_counter == 187)
	  estimate[338] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[338] <=  estimate[338];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[337] <= 0;
	else if(r_state == zStateEstimate & r_counter == 190)
	  estimate[337] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[337] <=  estimate[337];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[336] <= 0;
	else if(r_state == zStateEstimate & r_counter == 193)
	  estimate[336] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[336] <=  estimate[336];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[335] <= 0;
	else if(r_state == zStateEstimate & r_counter == 196)
	  estimate[335] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[335] <=  estimate[335];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[334] <= 0;
	else if(r_state == zStateEstimate & r_counter == 199)
	  estimate[334] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[334] <=  estimate[334];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[333] <= 0;
	else if(r_state == zStateEstimate & r_counter == 202)
	  estimate[333] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[333] <=  estimate[333];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[332] <= 0;
	else if(r_state == zStateEstimate & r_counter == 205)
	  estimate[332] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[332] <=  estimate[332];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[331] <= 0;
	else if(r_state == zStateEstimate & r_counter == 208)
	  estimate[331] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[331] <=  estimate[331];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[330] <= 0;
	else if(r_state == zStateEstimate & r_counter == 211)
	  estimate[330] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[330] <=  estimate[330];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[329] <= 0;
	else if(r_state == zStateEstimate & r_counter == 214)
	  estimate[329] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[329] <=  estimate[329];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[328] <= 0;
	else if(r_state == zStateEstimate & r_counter == 217)
	  estimate[328] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[328] <=  estimate[328];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[327] <= 0;
	else if(r_state == zStateEstimate & r_counter == 220)
	  estimate[327] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[327] <=  estimate[327];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[326] <= 0;
	else if(r_state == zStateEstimate & r_counter == 223)
	  estimate[326] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[326] <=  estimate[326];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[325] <= 0;
	else if(r_state == zStateEstimate & r_counter == 226)
	  estimate[325] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[325] <=  estimate[325];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[324] <= 0;
	else if(r_state == zStateEstimate & r_counter == 229)
	  estimate[324] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[324] <=  estimate[324];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[323] <= 0;
	else if(r_state == zStateEstimate & r_counter == 232)
	  estimate[323] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[323] <=  estimate[323];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[322] <= 0;
	else if(r_state == zStateEstimate & r_counter == 235)
	  estimate[322] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[322] <=  estimate[322];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[321] <= 0;
	else if(r_state == zStateEstimate & r_counter == 238)
	  estimate[321] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[321] <=  estimate[321];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[320] <= 0;
	else if(r_state == zStateEstimate & r_counter == 241)
	  estimate[320] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[320] <=  estimate[320];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[319] <= 0;
	else if(r_state == zStateEstimate & r_counter == 244)
	  estimate[319] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[319] <=  estimate[319];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[318] <= 0;
	else if(r_state == zStateEstimate & r_counter == 247)
	  estimate[318] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[318] <=  estimate[318];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[317] <= 0;
	else if(r_state == zStateEstimate & r_counter == 250)
	  estimate[317] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[317] <=  estimate[317];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[316] <= 0;
	else if(r_state == zStateEstimate & r_counter == 253)
	  estimate[316] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[316] <=  estimate[316];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[315] <= 0;
	else if(r_state == zStateEstimate & r_counter == 256)
	  estimate[315] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[315] <=  estimate[315];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[314] <= 0;
	else if(r_state == zStateEstimate & r_counter == 259)
	  estimate[314] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[314] <=  estimate[314];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[313] <= 0;
	else if(r_state == zStateEstimate & r_counter == 262)
	  estimate[313] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[313] <=  estimate[313];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[312] <= 0;
	else if(r_state == zStateEstimate & r_counter == 265)
	  estimate[312] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[312] <=  estimate[312];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[311] <= 0;
	else if(r_state == zStateEstimate & r_counter == 268)
	  estimate[311] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[311] <=  estimate[311];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[310] <= 0;
	else if(r_state == zStateEstimate & r_counter == 271)
	  estimate[310] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[310] <=  estimate[310];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[309] <= 0;
	else if(r_state == zStateEstimate & r_counter == 274)
	  estimate[309] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[309] <=  estimate[309];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[308] <= 0;
	else if(r_state == zStateEstimate & r_counter == 277)
	  estimate[308] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[308] <=  estimate[308];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[307] <= 0;
	else if(r_state == zStateEstimate & r_counter == 280)
	  estimate[307] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[307] <=  estimate[307];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[306] <= 0;
	else if(r_state == zStateEstimate & r_counter == 283)
	  estimate[306] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[306] <=  estimate[306];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[305] <= 0;
	else if(r_state == zStateEstimate & r_counter == 286)
	  estimate[305] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[305] <=  estimate[305];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[304] <= 0;
	else if(r_state == zStateEstimate & r_counter == 289)
	  estimate[304] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[304] <=  estimate[304];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[303] <= 0;
	else if(r_state == zStateEstimate & r_counter == 292)
	  estimate[303] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[303] <=  estimate[303];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[302] <= 0;
	else if(r_state == zStateEstimate & r_counter == 295)
	  estimate[302] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[302] <=  estimate[302];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[301] <= 0;
	else if(r_state == zStateEstimate & r_counter == 298)
	  estimate[301] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[301] <=  estimate[301];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[300] <= 0;
	else if(r_state == zStateEstimate & r_counter == 301)
	  estimate[300] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[300] <=  estimate[300];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[299] <= 0;
	else if(r_state == zStateEstimate & r_counter == 304)
	  estimate[299] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[299] <=  estimate[299];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[298] <= 0;
	else if(r_state == zStateEstimate & r_counter == 307)
	  estimate[298] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[298] <=  estimate[298];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[297] <= 0;
	else if(r_state == zStateEstimate & r_counter == 310)
	  estimate[297] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[297] <=  estimate[297];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[296] <= 0;
	else if(r_state == zStateEstimate & r_counter == 313)
	  estimate[296] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[296] <=  estimate[296];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[295] <= 0;
	else if(r_state == zStateEstimate & r_counter == 316)
	  estimate[295] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[295] <=  estimate[295];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[294] <= 0;
	else if(r_state == zStateEstimate & r_counter == 319)
	  estimate[294] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[294] <=  estimate[294];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[293] <= 0;
	else if(r_state == zStateEstimate & r_counter == 322)
	  estimate[293] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[293] <=  estimate[293];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[292] <= 0;
	else if(r_state == zStateEstimate & r_counter == 325)
	  estimate[292] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[292] <=  estimate[292];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[291] <= 0;
	else if(r_state == zStateEstimate & r_counter == 328)
	  estimate[291] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[291] <=  estimate[291];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[290] <= 0;
	else if(r_state == zStateEstimate & r_counter == 331)
	  estimate[290] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[290] <=  estimate[290];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[289] <= 0;
	else if(r_state == zStateEstimate & r_counter == 334)
	  estimate[289] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[289] <=  estimate[289];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[288] <= 0;
	else if(r_state == zStateEstimate & r_counter == 337)
	  estimate[288] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[288] <=  estimate[288];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[287] <= 0;
	else if(r_state == zStateEstimate & r_counter == 340)
	  estimate[287] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[287] <=  estimate[287];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[286] <= 0;
	else if(r_state == zStateEstimate & r_counter == 343)
	  estimate[286] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[286] <=  estimate[286];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[285] <= 0;
	else if(r_state == zStateEstimate & r_counter == 346)
	  estimate[285] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[285] <=  estimate[285];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[284] <= 0;
	else if(r_state == zStateEstimate & r_counter == 349)
	  estimate[284] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[284] <=  estimate[284];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[283] <= 0;
	else if(r_state == zStateEstimate & r_counter == 352)
	  estimate[283] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[283] <=  estimate[283];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[282] <= 0;
	else if(r_state == zStateEstimate & r_counter == 355)
	  estimate[282] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[282] <=  estimate[282];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[281] <= 0;
	else if(r_state == zStateEstimate & r_counter == 358)
	  estimate[281] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[281] <=  estimate[281];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[280] <= 0;
	else if(r_state == zStateEstimate & r_counter == 361)
	  estimate[280] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[280] <=  estimate[280];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[279] <= 0;
	else if(r_state == zStateEstimate & r_counter == 364)
	  estimate[279] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[279] <=  estimate[279];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[278] <= 0;
	else if(r_state == zStateEstimate & r_counter == 367)
	  estimate[278] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[278] <=  estimate[278];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[277] <= 0;
	else if(r_state == zStateEstimate & r_counter == 370)
	  estimate[277] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[277] <=  estimate[277];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[276] <= 0;
	else if(r_state == zStateEstimate & r_counter == 373)
	  estimate[276] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[276] <=  estimate[276];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[275] <= 0;
	else if(r_state == zStateEstimate & r_counter == 376)
	  estimate[275] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[275] <=  estimate[275];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[274] <= 0;
	else if(r_state == zStateEstimate & r_counter == 379)
	  estimate[274] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[274] <=  estimate[274];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[273] <= 0;
	else if(r_state == zStateEstimate & r_counter == 382)
	  estimate[273] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[273] <=  estimate[273];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[272] <= 0;
	else if(r_state == zStateEstimate & r_counter == 385)
	  estimate[272] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[272] <=  estimate[272];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[271] <= 0;
	else if(r_state == zStateEstimate & r_counter == 388)
	  estimate[271] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[271] <=  estimate[271];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[270] <= 0;
	else if(r_state == zStateEstimate & r_counter == 391)
	  estimate[270] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[270] <=  estimate[270];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[269] <= 0;
	else if(r_state == zStateEstimate & r_counter == 394)
	  estimate[269] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[269] <=  estimate[269];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[268] <= 0;
	else if(r_state == zStateEstimate & r_counter == 397)
	  estimate[268] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[268] <=  estimate[268];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[267] <= 0;
	else if(r_state == zStateEstimate & r_counter == 400)
	  estimate[267] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[267] <=  estimate[267];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[266] <= 0;
	else if(r_state == zStateEstimate & r_counter == 403)
	  estimate[266] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[266] <=  estimate[266];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[265] <= 0;
	else if(r_state == zStateEstimate & r_counter == 406)
	  estimate[265] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[265] <=  estimate[265];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[264] <= 0;
	else if(r_state == zStateEstimate & r_counter == 409)
	  estimate[264] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[264] <=  estimate[264];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[263] <= 0;
	else if(r_state == zStateEstimate & r_counter == 412)
	  estimate[263] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[263] <=  estimate[263];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[262] <= 0;
	else if(r_state == zStateEstimate & r_counter == 415)
	  estimate[262] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[262] <=  estimate[262];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[261] <= 0;
	else if(r_state == zStateEstimate & r_counter == 418)
	  estimate[261] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[261] <=  estimate[261];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[260] <= 0;
	else if(r_state == zStateEstimate & r_counter == 421)
	  estimate[260] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[260] <=  estimate[260];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[259] <= 0;
	else if(r_state == zStateEstimate & r_counter == 424)
	  estimate[259] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[259] <=  estimate[259];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[258] <= 0;
	else if(r_state == zStateEstimate & r_counter == 427)
	  estimate[258] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[258] <=  estimate[258];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[257] <= 0;
	else if(r_state == zStateEstimate & r_counter == 430)
	  estimate[257] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[257] <=  estimate[257];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[256] <= 0;
	else if(r_state == zStateEstimate & r_counter == 433)
	  estimate[256] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[256] <=  estimate[256];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[255] <= 0;
	else if(r_state == zStateEstimate & r_counter == 436)
	  estimate[255] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[255] <=  estimate[255];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[254] <= 0;
	else if(r_state == zStateEstimate & r_counter == 439)
	  estimate[254] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[254] <=  estimate[254];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[253] <= 0;
	else if(r_state == zStateEstimate & r_counter == 442)
	  estimate[253] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[253] <=  estimate[253];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[252] <= 0;
	else if(r_state == zStateEstimate & r_counter == 445)
	  estimate[252] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[252] <=  estimate[252];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[251] <= 0;
	else if(r_state == zStateEstimate & r_counter == 448)
	  estimate[251] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[251] <=  estimate[251];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[250] <= 0;
	else if(r_state == zStateEstimate & r_counter == 451)
	  estimate[250] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[250] <=  estimate[250];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[249] <= 0;
	else if(r_state == zStateEstimate & r_counter == 454)
	  estimate[249] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[249] <=  estimate[249];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[248] <= 0;
	else if(r_state == zStateEstimate & r_counter == 457)
	  estimate[248] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[248] <=  estimate[248];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[247] <= 0;
	else if(r_state == zStateEstimate & r_counter == 460)
	  estimate[247] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[247] <=  estimate[247];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[246] <= 0;
	else if(r_state == zStateEstimate & r_counter == 463)
	  estimate[246] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[246] <=  estimate[246];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[245] <= 0;
	else if(r_state == zStateEstimate & r_counter == 466)
	  estimate[245] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[245] <=  estimate[245];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[244] <= 0;
	else if(r_state == zStateEstimate & r_counter == 469)
	  estimate[244] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[244] <=  estimate[244];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[243] <= 0;
	else if(r_state == zStateEstimate & r_counter == 472)
	  estimate[243] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[243] <=  estimate[243];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[242] <= 0;
	else if(r_state == zStateEstimate & r_counter == 475)
	  estimate[242] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[242] <=  estimate[242];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[241] <= 0;
	else if(r_state == zStateEstimate & r_counter == 478)
	  estimate[241] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[241] <=  estimate[241];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[240] <= 0;
	else if(r_state == zStateEstimate & r_counter == 481)
	  estimate[240] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[240] <=  estimate[240];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[239] <= 0;
	else if(r_state == zStateEstimate & r_counter == 484)
	  estimate[239] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[239] <=  estimate[239];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[238] <= 0;
	else if(r_state == zStateEstimate & r_counter == 487)
	  estimate[238] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[238] <=  estimate[238];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[237] <= 0;
	else if(r_state == zStateEstimate & r_counter == 490)
	  estimate[237] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[237] <=  estimate[237];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[236] <= 0;
	else if(r_state == zStateEstimate & r_counter == 493)
	  estimate[236] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[236] <=  estimate[236];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[235] <= 0;
	else if(r_state == zStateEstimate & r_counter == 496)
	  estimate[235] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[235] <=  estimate[235];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[234] <= 0;
	else if(r_state == zStateEstimate & r_counter == 499)
	  estimate[234] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[234] <=  estimate[234];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[233] <= 0;
	else if(r_state == zStateEstimate & r_counter == 502)
	  estimate[233] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[233] <=  estimate[233];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[232] <= 0;
	else if(r_state == zStateEstimate & r_counter == 505)
	  estimate[232] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[232] <=  estimate[232];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[231] <= 0;
	else if(r_state == zStateEstimate & r_counter == 508)
	  estimate[231] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[231] <=  estimate[231];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[230] <= 0;
	else if(r_state == zStateEstimate & r_counter == 511)
	  estimate[230] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[230] <=  estimate[230];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[229] <= 0;
	else if(r_state == zStateEstimate & r_counter == 514)
	  estimate[229] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[229] <=  estimate[229];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[228] <= 0;
	else if(r_state == zStateEstimate & r_counter == 517)
	  estimate[228] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[228] <=  estimate[228];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[227] <= 0;
	else if(r_state == zStateEstimate & r_counter == 520)
	  estimate[227] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[227] <=  estimate[227];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[226] <= 0;
	else if(r_state == zStateEstimate & r_counter == 523)
	  estimate[226] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[226] <=  estimate[226];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[225] <= 0;
	else if(r_state == zStateEstimate & r_counter == 526)
	  estimate[225] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[225] <=  estimate[225];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[224] <= 0;
	else if(r_state == zStateEstimate & r_counter == 529)
	  estimate[224] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[224] <=  estimate[224];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[223] <= 0;
	else if(r_state == zStateEstimate & r_counter == 532)
	  estimate[223] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[223] <=  estimate[223];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[222] <= 0;
	else if(r_state == zStateEstimate & r_counter == 535)
	  estimate[222] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[222] <=  estimate[222];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[221] <= 0;
	else if(r_state == zStateEstimate & r_counter == 538)
	  estimate[221] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[221] <=  estimate[221];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[220] <= 0;
	else if(r_state == zStateEstimate & r_counter == 541)
	  estimate[220] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[220] <=  estimate[220];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[219] <= 0;
	else if(r_state == zStateEstimate & r_counter == 544)
	  estimate[219] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[219] <=  estimate[219];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[218] <= 0;
	else if(r_state == zStateEstimate & r_counter == 547)
	  estimate[218] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[218] <=  estimate[218];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[217] <= 0;
	else if(r_state == zStateEstimate & r_counter == 550)
	  estimate[217] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[217] <=  estimate[217];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[216] <= 0;
	else if(r_state == zStateEstimate & r_counter == 553)
	  estimate[216] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[216] <=  estimate[216];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[215] <= 0;
	else if(r_state == zStateEstimate & r_counter == 556)
	  estimate[215] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[215] <=  estimate[215];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[214] <= 0;
	else if(r_state == zStateEstimate & r_counter == 559)
	  estimate[214] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[214] <=  estimate[214];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[213] <= 0;
	else if(r_state == zStateEstimate & r_counter == 562)
	  estimate[213] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[213] <=  estimate[213];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[212] <= 0;
	else if(r_state == zStateEstimate & r_counter == 565)
	  estimate[212] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[212] <=  estimate[212];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[211] <= 0;
	else if(r_state == zStateEstimate & r_counter == 568)
	  estimate[211] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[211] <=  estimate[211];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[210] <= 0;
	else if(r_state == zStateEstimate & r_counter == 571)
	  estimate[210] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[210] <=  estimate[210];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[209] <= 0;
	else if(r_state == zStateEstimate & r_counter == 574)
	  estimate[209] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[209] <=  estimate[209];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[208] <= 0;
	else if(r_state == zStateEstimate & r_counter == 577)
	  estimate[208] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[208] <=  estimate[208];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[207] <= 0;
	else if(r_state == zStateEstimate & r_counter == 580)
	  estimate[207] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[207] <=  estimate[207];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[206] <= 0;
	else if(r_state == zStateEstimate & r_counter == 583)
	  estimate[206] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[206] <=  estimate[206];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[205] <= 0;
	else if(r_state == zStateEstimate & r_counter == 586)
	  estimate[205] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[205] <=  estimate[205];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[204] <= 0;
	else if(r_state == zStateEstimate & r_counter == 589)
	  estimate[204] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[204] <=  estimate[204];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[203] <= 0;
	else if(r_state == zStateEstimate & r_counter == 592)
	  estimate[203] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[203] <=  estimate[203];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[202] <= 0;
	else if(r_state == zStateEstimate & r_counter == 595)
	  estimate[202] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[202] <=  estimate[202];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[201] <= 0;
	else if(r_state == zStateEstimate & r_counter == 598)
	  estimate[201] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[201] <=  estimate[201];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[200] <= 0;
	else if(r_state == zStateEstimate & r_counter == 601)
	  estimate[200] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[200] <=  estimate[200];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[199] <= 0;
	else if(r_state == zStateEstimate & r_counter == 604)
	  estimate[199] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[199] <=  estimate[199];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[198] <= 0;
	else if(r_state == zStateEstimate & r_counter == 607)
	  estimate[198] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[198] <=  estimate[198];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[197] <= 0;
	else if(r_state == zStateEstimate & r_counter == 610)
	  estimate[197] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[197] <=  estimate[197];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[196] <= 0;
	else if(r_state == zStateEstimate & r_counter == 613)
	  estimate[196] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[196] <=  estimate[196];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[195] <= 0;
	else if(r_state == zStateEstimate & r_counter == 616)
	  estimate[195] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[195] <=  estimate[195];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[194] <= 0;
	else if(r_state == zStateEstimate & r_counter == 619)
	  estimate[194] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[194] <=  estimate[194];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[193] <= 0;
	else if(r_state == zStateEstimate & r_counter == 622)
	  estimate[193] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[193] <=  estimate[193];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[192] <= 0;
	else if(r_state == zStateEstimate & r_counter == 625)
	  estimate[192] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[192] <=  estimate[192];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[191] <= 0;
	else if(r_state == zStateEstimate & r_counter == 628)
	  estimate[191] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[191] <=  estimate[191];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[190] <= 0;
	else if(r_state == zStateEstimate & r_counter == 631)
	  estimate[190] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[190] <=  estimate[190];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[189] <= 0;
	else if(r_state == zStateEstimate & r_counter == 634)
	  estimate[189] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[189] <=  estimate[189];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[188] <= 0;
	else if(r_state == zStateEstimate & r_counter == 637)
	  estimate[188] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[188] <=  estimate[188];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[187] <= 0;
	else if(r_state == zStateEstimate & r_counter == 640)
	  estimate[187] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[187] <=  estimate[187];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[186] <= 0;
	else if(r_state == zStateEstimate & r_counter == 643)
	  estimate[186] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[186] <=  estimate[186];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[185] <= 0;
	else if(r_state == zStateEstimate & r_counter == 646)
	  estimate[185] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[185] <=  estimate[185];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[184] <= 0;
	else if(r_state == zStateEstimate & r_counter == 649)
	  estimate[184] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[184] <=  estimate[184];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[183] <= 0;
	else if(r_state == zStateEstimate & r_counter == 652)
	  estimate[183] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[183] <=  estimate[183];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[182] <= 0;
	else if(r_state == zStateEstimate & r_counter == 655)
	  estimate[182] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[182] <=  estimate[182];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[181] <= 0;
	else if(r_state == zStateEstimate & r_counter == 658)
	  estimate[181] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[181] <=  estimate[181];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[180] <= 0;
	else if(r_state == zStateEstimate & r_counter == 661)
	  estimate[180] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[180] <=  estimate[180];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[179] <= 0;
	else if(r_state == zStateEstimate & r_counter == 664)
	  estimate[179] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[179] <=  estimate[179];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[178] <= 0;
	else if(r_state == zStateEstimate & r_counter == 667)
	  estimate[178] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[178] <=  estimate[178];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[177] <= 0;
	else if(r_state == zStateEstimate & r_counter == 670)
	  estimate[177] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[177] <=  estimate[177];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[176] <= 0;
	else if(r_state == zStateEstimate & r_counter == 673)
	  estimate[176] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[176] <=  estimate[176];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[175] <= 0;
	else if(r_state == zStateEstimate & r_counter == 676)
	  estimate[175] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[175] <=  estimate[175];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[174] <= 0;
	else if(r_state == zStateEstimate & r_counter == 679)
	  estimate[174] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[174] <=  estimate[174];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[173] <= 0;
	else if(r_state == zStateEstimate & r_counter == 682)
	  estimate[173] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[173] <=  estimate[173];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[172] <= 0;
	else if(r_state == zStateEstimate & r_counter == 685)
	  estimate[172] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[172] <=  estimate[172];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[171] <= 0;
	else if(r_state == zStateEstimate & r_counter == 688)
	  estimate[171] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[171] <=  estimate[171];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[170] <= 0;
	else if(r_state == zStateEstimate & r_counter == 691)
	  estimate[170] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[170] <=  estimate[170];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[169] <= 0;
	else if(r_state == zStateEstimate & r_counter == 694)
	  estimate[169] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[169] <=  estimate[169];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[168] <= 0;
	else if(r_state == zStateEstimate & r_counter == 697)
	  estimate[168] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[168] <=  estimate[168];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[167] <= 0;
	else if(r_state == zStateEstimate & r_counter == 700)
	  estimate[167] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[167] <=  estimate[167];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[166] <= 0;
	else if(r_state == zStateEstimate & r_counter == 703)
	  estimate[166] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[166] <=  estimate[166];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[165] <= 0;
	else if(r_state == zStateEstimate & r_counter == 706)
	  estimate[165] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[165] <=  estimate[165];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[164] <= 0;
	else if(r_state == zStateEstimate & r_counter == 709)
	  estimate[164] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[164] <=  estimate[164];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[163] <= 0;
	else if(r_state == zStateEstimate & r_counter == 712)
	  estimate[163] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[163] <=  estimate[163];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[162] <= 0;
	else if(r_state == zStateEstimate & r_counter == 715)
	  estimate[162] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[162] <=  estimate[162];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[161] <= 0;
	else if(r_state == zStateEstimate & r_counter == 718)
	  estimate[161] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[161] <=  estimate[161];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[160] <= 0;
	else if(r_state == zStateEstimate & r_counter == 721)
	  estimate[160] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[160] <=  estimate[160];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[159] <= 0;
	else if(r_state == zStateEstimate & r_counter == 724)
	  estimate[159] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[159] <=  estimate[159];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[158] <= 0;
	else if(r_state == zStateEstimate & r_counter == 727)
	  estimate[158] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[158] <=  estimate[158];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[157] <= 0;
	else if(r_state == zStateEstimate & r_counter == 730)
	  estimate[157] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[157] <=  estimate[157];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[156] <= 0;
	else if(r_state == zStateEstimate & r_counter == 733)
	  estimate[156] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[156] <=  estimate[156];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[155] <= 0;
	else if(r_state == zStateEstimate & r_counter == 736)
	  estimate[155] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[155] <=  estimate[155];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[154] <= 0;
	else if(r_state == zStateEstimate & r_counter == 739)
	  estimate[154] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[154] <=  estimate[154];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[153] <= 0;
	else if(r_state == zStateEstimate & r_counter == 742)
	  estimate[153] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[153] <=  estimate[153];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[152] <= 0;
	else if(r_state == zStateEstimate & r_counter == 745)
	  estimate[152] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[152] <=  estimate[152];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[151] <= 0;
	else if(r_state == zStateEstimate & r_counter == 748)
	  estimate[151] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[151] <=  estimate[151];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[150] <= 0;
	else if(r_state == zStateEstimate & r_counter == 751)
	  estimate[150] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[150] <=  estimate[150];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[149] <= 0;
	else if(r_state == zStateEstimate & r_counter == 754)
	  estimate[149] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[149] <=  estimate[149];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[148] <= 0;
	else if(r_state == zStateEstimate & r_counter == 757)
	  estimate[148] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[148] <=  estimate[148];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[147] <= 0;
	else if(r_state == zStateEstimate & r_counter == 760)
	  estimate[147] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[147] <=  estimate[147];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[146] <= 0;
	else if(r_state == zStateEstimate & r_counter == 763)
	  estimate[146] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[146] <=  estimate[146];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[145] <= 0;
	else if(r_state == zStateEstimate & r_counter == 766)
	  estimate[145] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[145] <=  estimate[145];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[144] <= 0;
	else if(r_state == zStateEstimate & r_counter == 769)
	  estimate[144] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[144] <=  estimate[144];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[143] <= 0;
	else if(r_state == zStateEstimate & r_counter == 772)
	  estimate[143] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[143] <=  estimate[143];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[142] <= 0;
	else if(r_state == zStateEstimate & r_counter == 775)
	  estimate[142] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[142] <=  estimate[142];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[141] <= 0;
	else if(r_state == zStateEstimate & r_counter == 778)
	  estimate[141] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[141] <=  estimate[141];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[140] <= 0;
	else if(r_state == zStateEstimate & r_counter == 781)
	  estimate[140] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[140] <=  estimate[140];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[139] <= 0;
	else if(r_state == zStateEstimate & r_counter == 784)
	  estimate[139] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[139] <=  estimate[139];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[138] <= 0;
	else if(r_state == zStateEstimate & r_counter == 787)
	  estimate[138] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[138] <=  estimate[138];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[137] <= 0;
	else if(r_state == zStateEstimate & r_counter == 790)
	  estimate[137] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[137] <=  estimate[137];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[136] <= 0;
	else if(r_state == zStateEstimate & r_counter == 793)
	  estimate[136] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[136] <=  estimate[136];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[135] <= 0;
	else if(r_state == zStateEstimate & r_counter == 796)
	  estimate[135] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[135] <=  estimate[135];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[134] <= 0;
	else if(r_state == zStateEstimate & r_counter == 799)
	  estimate[134] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[134] <=  estimate[134];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[133] <= 0;
	else if(r_state == zStateEstimate & r_counter == 802)
	  estimate[133] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[133] <=  estimate[133];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[132] <= 0;
	else if(r_state == zStateEstimate & r_counter == 805)
	  estimate[132] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[132] <=  estimate[132];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[131] <= 0;
	else if(r_state == zStateEstimate & r_counter == 808)
	  estimate[131] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[131] <=  estimate[131];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[130] <= 0;
	else if(r_state == zStateEstimate & r_counter == 811)
	  estimate[130] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[130] <=  estimate[130];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[129] <= 0;
	else if(r_state == zStateEstimate & r_counter == 814)
	  estimate[129] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[129] <=  estimate[129];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[128] <= 0;
	else if(r_state == zStateEstimate & r_counter == 817)
	  estimate[128] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[128] <=  estimate[128];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[127] <= 0;
	else if(r_state == zStateEstimate & r_counter == 820)
	  estimate[127] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[127] <=  estimate[127];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[126] <= 0;
	else if(r_state == zStateEstimate & r_counter == 823)
	  estimate[126] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[126] <=  estimate[126];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[125] <= 0;
	else if(r_state == zStateEstimate & r_counter == 826)
	  estimate[125] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[125] <=  estimate[125];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[124] <= 0;
	else if(r_state == zStateEstimate & r_counter == 829)
	  estimate[124] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[124] <=  estimate[124];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[123] <= 0;
	else if(r_state == zStateEstimate & r_counter == 832)
	  estimate[123] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[123] <=  estimate[123];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[122] <= 0;
	else if(r_state == zStateEstimate & r_counter == 835)
	  estimate[122] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[122] <=  estimate[122];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[121] <= 0;
	else if(r_state == zStateEstimate & r_counter == 838)
	  estimate[121] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[121] <=  estimate[121];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[120] <= 0;
	else if(r_state == zStateEstimate & r_counter == 841)
	  estimate[120] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[120] <=  estimate[120];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[119] <= 0;
	else if(r_state == zStateEstimate & r_counter == 844)
	  estimate[119] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[119] <=  estimate[119];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[118] <= 0;
	else if(r_state == zStateEstimate & r_counter == 847)
	  estimate[118] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[118] <=  estimate[118];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[117] <= 0;
	else if(r_state == zStateEstimate & r_counter == 850)
	  estimate[117] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[117] <=  estimate[117];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[116] <= 0;
	else if(r_state == zStateEstimate & r_counter == 853)
	  estimate[116] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[116] <=  estimate[116];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[115] <= 0;
	else if(r_state == zStateEstimate & r_counter == 856)
	  estimate[115] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[115] <=  estimate[115];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[114] <= 0;
	else if(r_state == zStateEstimate & r_counter == 859)
	  estimate[114] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[114] <=  estimate[114];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[113] <= 0;
	else if(r_state == zStateEstimate & r_counter == 862)
	  estimate[113] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[113] <=  estimate[113];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[112] <= 0;
	else if(r_state == zStateEstimate & r_counter == 865)
	  estimate[112] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[112] <=  estimate[112];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[111] <= 0;
	else if(r_state == zStateEstimate & r_counter == 868)
	  estimate[111] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[111] <=  estimate[111];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[110] <= 0;
	else if(r_state == zStateEstimate & r_counter == 871)
	  estimate[110] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[110] <=  estimate[110];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[109] <= 0;
	else if(r_state == zStateEstimate & r_counter == 874)
	  estimate[109] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[109] <=  estimate[109];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[108] <= 0;
	else if(r_state == zStateEstimate & r_counter == 877)
	  estimate[108] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[108] <=  estimate[108];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[107] <= 0;
	else if(r_state == zStateEstimate & r_counter == 880)
	  estimate[107] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[107] <=  estimate[107];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[106] <= 0;
	else if(r_state == zStateEstimate & r_counter == 883)
	  estimate[106] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[106] <=  estimate[106];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[105] <= 0;
	else if(r_state == zStateEstimate & r_counter == 886)
	  estimate[105] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[105] <=  estimate[105];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[104] <= 0;
	else if(r_state == zStateEstimate & r_counter == 889)
	  estimate[104] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[104] <=  estimate[104];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[103] <= 0;
	else if(r_state == zStateEstimate & r_counter == 892)
	  estimate[103] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[103] <=  estimate[103];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[102] <= 0;
	else if(r_state == zStateEstimate & r_counter == 895)
	  estimate[102] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[102] <=  estimate[102];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[101] <= 0;
	else if(r_state == zStateEstimate & r_counter == 898)
	  estimate[101] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[101] <=  estimate[101];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[100] <= 0;
	else if(r_state == zStateEstimate & r_counter == 901)
	  estimate[100] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[100] <=  estimate[100];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[99] <= 0;
	else if(r_state == zStateEstimate & r_counter == 904)
	  estimate[99] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[99] <=  estimate[99];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[98] <= 0;
	else if(r_state == zStateEstimate & r_counter == 907)
	  estimate[98] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[98] <=  estimate[98];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[97] <= 0;
	else if(r_state == zStateEstimate & r_counter == 910)
	  estimate[97] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[97] <=  estimate[97];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[96] <= 0;
	else if(r_state == zStateEstimate & r_counter == 913)
	  estimate[96] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[96] <=  estimate[96];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[95] <= 0;
	else if(r_state == zStateEstimate & r_counter == 916)
	  estimate[95] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[95] <=  estimate[95];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[94] <= 0;
	else if(r_state == zStateEstimate & r_counter == 919)
	  estimate[94] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[94] <=  estimate[94];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[93] <= 0;
	else if(r_state == zStateEstimate & r_counter == 922)
	  estimate[93] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[93] <=  estimate[93];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[92] <= 0;
	else if(r_state == zStateEstimate & r_counter == 925)
	  estimate[92] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[92] <=  estimate[92];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[91] <= 0;
	else if(r_state == zStateEstimate & r_counter == 928)
	  estimate[91] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[91] <=  estimate[91];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[90] <= 0;
	else if(r_state == zStateEstimate & r_counter == 931)
	  estimate[90] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[90] <=  estimate[90];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[89] <= 0;
	else if(r_state == zStateEstimate & r_counter == 934)
	  estimate[89] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[89] <=  estimate[89];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[88] <= 0;
	else if(r_state == zStateEstimate & r_counter == 937)
	  estimate[88] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[88] <=  estimate[88];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[87] <= 0;
	else if(r_state == zStateEstimate & r_counter == 940)
	  estimate[87] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[87] <=  estimate[87];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[86] <= 0;
	else if(r_state == zStateEstimate & r_counter == 943)
	  estimate[86] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[86] <=  estimate[86];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[85] <= 0;
	else if(r_state == zStateEstimate & r_counter == 946)
	  estimate[85] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[85] <=  estimate[85];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[84] <= 0;
	else if(r_state == zStateEstimate & r_counter == 949)
	  estimate[84] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[84] <=  estimate[84];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[83] <= 0;
	else if(r_state == zStateEstimate & r_counter == 952)
	  estimate[83] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[83] <=  estimate[83];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[82] <= 0;
	else if(r_state == zStateEstimate & r_counter == 955)
	  estimate[82] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[82] <=  estimate[82];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[81] <= 0;
	else if(r_state == zStateEstimate & r_counter == 958)
	  estimate[81] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[81] <=  estimate[81];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[80] <= 0;
	else if(r_state == zStateEstimate & r_counter == 961)
	  estimate[80] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[80] <=  estimate[80];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[79] <= 0;
	else if(r_state == zStateEstimate & r_counter == 964)
	  estimate[79] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[79] <=  estimate[79];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[78] <= 0;
	else if(r_state == zStateEstimate & r_counter == 967)
	  estimate[78] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[78] <=  estimate[78];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[77] <= 0;
	else if(r_state == zStateEstimate & r_counter == 970)
	  estimate[77] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[77] <=  estimate[77];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[76] <= 0;
	else if(r_state == zStateEstimate & r_counter == 973)
	  estimate[76] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[76] <=  estimate[76];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[75] <= 0;
	else if(r_state == zStateEstimate & r_counter == 976)
	  estimate[75] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[75] <=  estimate[75];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[74] <= 0;
	else if(r_state == zStateEstimate & r_counter == 979)
	  estimate[74] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[74] <=  estimate[74];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[73] <= 0;
	else if(r_state == zStateEstimate & r_counter == 982)
	  estimate[73] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[73] <=  estimate[73];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[72] <= 0;
	else if(r_state == zStateEstimate & r_counter == 985)
	  estimate[72] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[72] <=  estimate[72];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[71] <= 0;
	else if(r_state == zStateEstimate & r_counter == 988)
	  estimate[71] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[71] <=  estimate[71];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[70] <= 0;
	else if(r_state == zStateEstimate & r_counter == 991)
	  estimate[70] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[70] <=  estimate[70];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[69] <= 0;
	else if(r_state == zStateEstimate & r_counter == 994)
	  estimate[69] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[69] <=  estimate[69];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[68] <= 0;
	else if(r_state == zStateEstimate & r_counter == 997)
	  estimate[68] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[68] <=  estimate[68];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[67] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1000)
	  estimate[67] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[67] <=  estimate[67];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[66] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1003)
	  estimate[66] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[66] <=  estimate[66];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[65] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1006)
	  estimate[65] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[65] <=  estimate[65];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[64] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1009)
	  estimate[64] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[64] <=  estimate[64];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[63] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1012)
	  estimate[63] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[63] <=  estimate[63];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[62] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1015)
	  estimate[62] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[62] <=  estimate[62];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[61] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1018)
	  estimate[61] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[61] <=  estimate[61];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[60] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1021)
	  estimate[60] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[60] <=  estimate[60];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[59] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1024)
	  estimate[59] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[59] <=  estimate[59];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[58] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1027)
	  estimate[58] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[58] <=  estimate[58];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[57] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1030)
	  estimate[57] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[57] <=  estimate[57];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[56] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1033)
	  estimate[56] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[56] <=  estimate[56];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[55] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1036)
	  estimate[55] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[55] <=  estimate[55];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[54] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1039)
	  estimate[54] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[54] <=  estimate[54];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[53] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1042)
	  estimate[53] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[53] <=  estimate[53];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[52] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1045)
	  estimate[52] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[52] <=  estimate[52];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[51] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1048)
	  estimate[51] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[51] <=  estimate[51];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[50] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1051)
	  estimate[50] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[50] <=  estimate[50];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[49] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1054)
	  estimate[49] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[49] <=  estimate[49];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[48] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1057)
	  estimate[48] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[48] <=  estimate[48];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[47] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1060)
	  estimate[47] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[47] <=  estimate[47];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[46] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1063)
	  estimate[46] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[46] <=  estimate[46];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[45] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1066)
	  estimate[45] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[45] <=  estimate[45];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[44] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1069)
	  estimate[44] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[44] <=  estimate[44];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[43] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1072)
	  estimate[43] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[43] <=  estimate[43];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[42] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1075)
	  estimate[42] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[42] <=  estimate[42];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[41] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1078)
	  estimate[41] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[41] <=  estimate[41];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[40] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1081)
	  estimate[40] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[40] <=  estimate[40];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[39] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1084)
	  estimate[39] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[39] <=  estimate[39];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[38] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1087)
	  estimate[38] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[38] <=  estimate[38];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[37] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1090)
	  estimate[37] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[37] <=  estimate[37];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[36] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1093)
	  estimate[36] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[36] <=  estimate[36];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[35] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1096)
	  estimate[35] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[35] <=  estimate[35];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[34] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1099)
	  estimate[34] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[34] <=  estimate[34];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[33] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1102)
	  estimate[33] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[33] <=  estimate[33];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[32] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1105)
	  estimate[32] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[32] <=  estimate[32];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[31] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1108)
	  estimate[31] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[31] <=  estimate[31];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[30] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1111)
	  estimate[30] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[30] <=  estimate[30];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[29] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1114)
	  estimate[29] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[29] <=  estimate[29];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[28] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1117)
	  estimate[28] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[28] <=  estimate[28];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[27] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1120)
	  estimate[27] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[27] <=  estimate[27];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[26] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1123)
	  estimate[26] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[26] <=  estimate[26];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[25] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1126)
	  estimate[25] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[25] <=  estimate[25];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[24] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1129)
	  estimate[24] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[24] <=  estimate[24];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[23] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1132)
	  estimate[23] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[23] <=  estimate[23];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[22] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1135)
	  estimate[22] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[22] <=  estimate[22];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[21] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1138)
	  estimate[21] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[21] <=  estimate[21];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[20] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1141)
	  estimate[20] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[20] <=  estimate[20];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[19] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1144)
	  estimate[19] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[19] <=  estimate[19];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[18] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1147)
	  estimate[18] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[18] <=  estimate[18];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[17] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1150)
	  estimate[17] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[17] <=  estimate[17];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[16] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1153)
	  estimate[16] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[16] <=  estimate[16];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[15] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1156)
	  estimate[15] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[15] <=  estimate[15];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[14] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1159)
	  estimate[14] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[14] <=  estimate[14];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[13] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1162)
	  estimate[13] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[13] <=  estimate[13];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[12] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1165)
	  estimate[12] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[12] <=  estimate[12];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[11] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1168)
	  estimate[11] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[11] <=  estimate[11];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[10] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1171)
	  estimate[10] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[10] <=  estimate[10];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[9] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1174)
	  estimate[9] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[9] <=  estimate[9];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[8] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1177)
	  estimate[8] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[8] <=  estimate[8];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[7] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1180)
	  estimate[7] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[7] <=  estimate[7];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[6] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1183)
	  estimate[6] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[6] <=  estimate[6];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[5] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1186)
	  estimate[5] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[5] <=  estimate[5];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[4] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1189)
	  estimate[4] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[4] <=  estimate[4];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[3] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1192)
	  estimate[3] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[3] <=  estimate[3];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[2] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1195)
	  estimate[2] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[2] <=  estimate[2];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[1] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1198)
	  estimate[1] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[1] <=  estimate[1];
     end
   /**/
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  estimate[0] <= 0;
	else if(r_state == zStateEstimate & r_counter == 1201)
	  estimate[0] <= (o_data_test_beta > 0) ? 0:1;
	else
	  estimate[0] <=  estimate[0];
     end
   /**/
	

   
   
   //行処理が終わった時にパリティビットが1であれば出力valid信号を1とする
   assign o_val = ( (r_state==zStateColumn) & (r_counter == 2) & (parity==1) ) ? 1:0;
   
   //sram関係

   //lambda
   assign i_wen_lambda=(r_state==zStateLambdaInit) ? 1:0;
   assign i_waddr_lambda=r_counter;
   assign i_raddr_lambda=/**/
			 (r_state == zStateBetaInit) & (r_counter == 0) ? 125:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 1) ? 201:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 2) ? 202:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 3) ? 203:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 4) ? 204:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 5) ? 205:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 6) ? 206:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 7) ? 207:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 8) ? 208:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 9) ? 209:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 10) ? 210:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 11) ? 211:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 12) ? 212:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 13) ? 213:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 14) ? 214:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 15) ? 215:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 16) ? 216:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 17) ? 217:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 18) ? 218:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 19) ? 219:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 20) ? 220:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 21) ? 221:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 22) ? 222:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 23) ? 223:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 24) ? 224:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 25) ? 225:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 26) ? 226:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 27) ? 227:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 28) ? 228:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 29) ? 229:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 30) ? 230:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 31) ? 231:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 32) ? 232:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 33) ? 233:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 34) ? 234:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 35) ? 235:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 36) ? 236:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 37) ? 237:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 38) ? 238:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 39) ? 239:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 40) ? 240:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 41) ? 241:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 42) ? 242:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 43) ? 243:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 44) ? 244:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 45) ? 245:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 46) ? 246:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 47) ? 247:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 48) ? 9:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 49) ? 248:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 50) ? 249:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 51) ? 250:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 52) ? 251:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 53) ? 252:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 54) ? 253:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 55) ? 254:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 56) ? 255:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 57) ? 256:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 58) ? 257:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 59) ? 258:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 60) ? 259:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 61) ? 260:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 62) ? 261:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 63) ? 262:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 64) ? 61:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 65) ? 263:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 66) ? 264:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 67) ? 265:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 68) ? 266:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 69) ? 267:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 70) ? 268:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 71) ? 269:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 72) ? 29:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 73) ? 270:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 74) ? 271:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 75) ? 272:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 76) ? 273:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 77) ? 274:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 78) ? 275:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 79) ? 276:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 80) ? 277:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 81) ? 278:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 82) ? 279:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 83) ? 280:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 84) ? 101:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 85) ? 281:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 86) ? 282:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 87) ? 283:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 88) ? 13:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 89) ? 284:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 90) ? 285:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 91) ? 286:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 92) ? 287:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 93) ? 288:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 94) ? 289:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 95) ? 290:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 96) ? 53:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 97) ? 54:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 98) ? 291:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 99) ? 292:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 100) ? 157:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 101) ? 293:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 102) ? 294:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 103) ? 295:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 104) ? 296:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 105) ? 297:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 106) ? 298:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 107) ? 299:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 108) ? 65:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 109) ? 300:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 110) ? 301:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 111) ? 302:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 112) ? 5:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 113) ? 173:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 114) ? 303:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 115) ? 304:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 116) ? 17:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 117) ? 21:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 118) ? 305:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 119) ? 306:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 120) ? 33:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 121) ? 41:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 122) ? 49:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 123) ? 307:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 124) ? 57:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 125) ? 308:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 126) ? 309:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 127) ? 310:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 128) ? 69:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 129) ? 85:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 130) ? 97:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 131) ? 311:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 132) ? 105:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 133) ? 110:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 134) ? 121:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 135) ? 312:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 136) ? 129:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 137) ? 133:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 138) ? 141:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 139) ? 313:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 140) ? 1:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 141) ? 189:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 142) ? 314:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 143) ? 315:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 144) ? 16:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 145) ? 316:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 146) ? 317:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 147) ? 318:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 148) ? 23:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 149) ? 25:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 150) ? 319:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 151) ? 320:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 152) ? 30:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 153) ? 37:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 154) ? 321:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 155) ? 322:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 156) ? 45:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 157) ? 323:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 158) ? 324:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 159) ? 325:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 160) ? 326:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 161) ? 327:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 162) ? 328:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 163) ? 329:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 164) ? 73:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 165) ? 77:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 166) ? 81:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 167) ? 330:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 168) ? 89:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 169) ? 91:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 170) ? 93:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 171) ? 331:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 172) ? 109:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 173) ? 332:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 174) ? 333:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 175) ? 334:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 176) ? 113:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 177) ? 117:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 178) ? 335:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 179) ? 336:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 180) ? 137:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 181) ? 337:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 182) ? 338:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 183) ? 339:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 184) ? 145:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 185) ? 149:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 186) ? 153:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 187) ? 340:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 188) ? 161:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 189) ? 165:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 190) ? 169:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 191) ? 341:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 192) ? 177:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 193) ? 181:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 194) ? 185:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 195) ? 342:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 196) ? 0:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 197) ? 193:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 198) ? 197:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 199) ? 343:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 200) ? 2:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 201) ? 3:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 202) ? 4:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 203) ? 344:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 204) ? 6:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 205) ? 7:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 206) ? 8:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 207) ? 345:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 208) ? 10:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 209) ? 11:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 210) ? 12:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 211) ? 346:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 212) ? 14:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 213) ? 15:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 214) ? 347:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 215) ? 348:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 216) ? 18:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 217) ? 19:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 218) ? 20:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 219) ? 349:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 220) ? 22:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 221) ? 24:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 222) ? 350:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 223) ? 351:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 224) ? 26:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 225) ? 27:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 226) ? 28:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 227) ? 352:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 228) ? 31:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 229) ? 32:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 230) ? 353:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 231) ? 354:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 232) ? 34:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 233) ? 35:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 234) ? 36:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 235) ? 355:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 236) ? 38:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 237) ? 39:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 238) ? 40:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 239) ? 356:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 240) ? 42:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 241) ? 43:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 242) ? 44:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 243) ? 357:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 244) ? 46:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 245) ? 47:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 246) ? 48:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 247) ? 358:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 248) ? 50:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 249) ? 51:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 250) ? 52:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 251) ? 359:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 252) ? 55:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 253) ? 56:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 254) ? 360:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 255) ? 361:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 256) ? 58:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 257) ? 59:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 258) ? 60:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 259) ? 362:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 260) ? 62:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 261) ? 63:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 262) ? 64:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 263) ? 363:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 264) ? 66:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 265) ? 67:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 266) ? 68:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 267) ? 364:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 268) ? 70:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 269) ? 71:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 270) ? 72:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 271) ? 365:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 272) ? 74:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 273) ? 75:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 274) ? 76:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 275) ? 366:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 276) ? 78:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 277) ? 79:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 278) ? 80:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 279) ? 367:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 280) ? 82:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 281) ? 83:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 282) ? 84:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 283) ? 368:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 284) ? 86:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 285) ? 87:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 286) ? 88:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 287) ? 369:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 288) ? 90:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 289) ? 92:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 290) ? 370:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 291) ? 371:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 292) ? 94:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 293) ? 95:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 294) ? 96:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 295) ? 372:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 296) ? 98:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 297) ? 99:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 298) ? 100:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 299) ? 373:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 300) ? 102:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 301) ? 103:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 302) ? 104:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 303) ? 374:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 304) ? 106:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 305) ? 107:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 306) ? 108:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 307) ? 375:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 308) ? 111:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 309) ? 112:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 310) ? 376:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 311) ? 377:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 312) ? 114:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 313) ? 115:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 314) ? 116:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 315) ? 378:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 316) ? 118:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 317) ? 119:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 318) ? 120:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 319) ? 379:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 320) ? 122:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 321) ? 123:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 322) ? 124:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 323) ? 380:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 324) ? 126:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 325) ? 127:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 326) ? 128:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 327) ? 381:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 328) ? 130:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 329) ? 131:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 330) ? 132:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 331) ? 382:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 332) ? 134:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 333) ? 135:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 334) ? 136:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 335) ? 383:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 336) ? 138:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 337) ? 139:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 338) ? 140:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 339) ? 384:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 340) ? 142:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 341) ? 143:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 342) ? 144:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 343) ? 385:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 344) ? 146:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 345) ? 147:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 346) ? 148:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 347) ? 386:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 348) ? 150:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 349) ? 151:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 350) ? 152:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 351) ? 387:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 352) ? 154:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 353) ? 155:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 354) ? 156:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 355) ? 388:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 356) ? 158:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 357) ? 159:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 358) ? 160:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 359) ? 389:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 360) ? 162:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 361) ? 163:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 362) ? 164:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 363) ? 390:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 364) ? 166:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 365) ? 167:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 366) ? 168:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 367) ? 391:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 368) ? 170:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 369) ? 171:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 370) ? 172:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 371) ? 392:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 372) ? 174:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 373) ? 175:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 374) ? 176:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 375) ? 393:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 376) ? 178:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 377) ? 179:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 378) ? 180:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 379) ? 394:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 380) ? 182:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 381) ? 183:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 382) ? 184:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 383) ? 395:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 384) ? 186:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 385) ? 187:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 386) ? 188:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 387) ? 396:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 388) ? 190:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 389) ? 191:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 390) ? 192:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 391) ? 397:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 392) ? 194:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 393) ? 195:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 394) ? 196:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 395) ? 398:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 396) ? 198:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 397) ? 199:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 398) ? 200:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 399) ? 399:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 400) ? 74:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 401) ? 135:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 402) ? 178:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 403) ? 325:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 404) ? 205:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 405) ? 236:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 406) ? 285:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 407) ? 335:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 408) ? 22:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 409) ? 82:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 410) ? 334:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 411) ? 391:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 412) ? 113:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 413) ? 126:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 414) ? 298:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 415) ? 329:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 416) ? 8:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 417) ? 69:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 418) ? 295:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 419) ? 385:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 420) ? 11:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 421) ? 198:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 422) ? 207:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 423) ? 332:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 424) ? 189:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 425) ? 258:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 426) ? 271:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 427) ? 346:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 428) ? 46:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 429) ? 65:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 430) ? 300:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 431) ? 347:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 432) ? 52:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 433) ? 101:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 434) ? 210:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 435) ? 376:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 436) ? 37:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 437) ? 110:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 438) ? 196:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 439) ? 257:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 440) ? 161:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 441) ? 277:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 442) ? 312:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 443) ? 356:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 444) ? 98:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 445) ? 112:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 446) ? 174:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 447) ? 317:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 448) ? 61:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 449) ? 88:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 450) ? 130:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 451) ? 250:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 452) ? 131:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 453) ? 199:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 454) ? 377:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 455) ? 399:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 456) ? 64:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 457) ? 102:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 458) ? 324:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 459) ? 368:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 460) ? 254:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 461) ? 343:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 462) ? 359:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 463) ? 372:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 464) ? 10:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 465) ? 30:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 466) ? 180:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 467) ? 243:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 468) ? 105:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 469) ? 228:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 470) ? 331:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 471) ? 365:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 472) ? 18:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 473) ? 79:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 474) ? 226:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 475) ? 296:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 476) ? 13:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 477) ? 150:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 478) ? 194:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 479) ? 280:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 480) ? 96:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 481) ? 136:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 482) ? 195:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 483) ? 315:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 484) ? 119:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 485) ? 129:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 486) ? 252:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 487) ? 353:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 488) ? 173:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 489) ? 202:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 490) ? 223:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 491) ? 389:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 492) ? 50:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 493) ? 137:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 494) ? 229:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 495) ? 272:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 496) ? 16:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 497) ? 40:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 498) ? 86:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 499) ? 293:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 500) ? 99:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 501) ? 221:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 502) ? 244:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 503) ? 267:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 504) ? 38:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 505) ? 95:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 506) ? 184:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 507) ? 327:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 508) ? 53:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 509) ? 206:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 510) ? 242:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 511) ? 248:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 512) ? 3:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 513) ? 72:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 514) ? 238:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 515) ? 383:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 516) ? 45:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 517) ? 212:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 518) ? 251:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 519) ? 379:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 520) ? 168:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 521) ? 182:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 522) ? 299:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 523) ? 392:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 524) ? 78:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 525) ? 190:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 526) ? 286:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 527) ? 384:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 528) ? 59:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 529) ? 67:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 530) ? 187:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 531) ? 354:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 532) ? 89:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 533) ? 108:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 534) ? 274:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 535) ? 375:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 536) ? 153:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 537) ? 213:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 538) ? 246:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 539) ? 398:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 540) ? 36:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 541) ? 261:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 542) ? 270:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 543) ? 283:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 544) ? 118:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 545) ? 144:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 546) ? 151:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 547) ? 371:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 548) ? 76:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 549) ? 107:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 550) ? 292:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 551) ? 330:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 552) ? 25:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 553) ? 35:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 554) ? 214:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 555) ? 294:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 556) ? 49:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 557) ? 162:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 558) ? 224:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 559) ? 382:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 560) ? 5:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 561) ? 209:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 562) ? 273:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 563) ? 344:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 564) ? 34:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 565) ? 125:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 566) ? 201:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 567) ? 319:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 568) ? 140:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 569) ? 146:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 570) ? 320:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 571) ? 388:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 572) ? 19:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 573) ? 183:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 574) ? 310:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 575) ? 373:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 576) ? 48:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 577) ? 57:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 578) ? 170:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 579) ? 234:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 580) ? 116:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 581) ? 239:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 582) ? 350:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 583) ? 364:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 584) ? 32:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 585) ? 127:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 586) ? 152:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 587) ? 328:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 588) ? 142:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 589) ? 188:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 590) ? 360:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 591) ? 396:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 592) ? 158:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 593) ? 218:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 594) ? 266:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 595) ? 352:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 596) ? 166:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 597) ? 249:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 598) ? 276:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 599) ? 323:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 600) ? 43:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 601) ? 197:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 602) ? 219:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 603) ? 290:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 604) ? 14:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 605) ? 231:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 606) ? 278:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 607) ? 387:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 608) ? 62:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 609) ? 122:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 610) ? 143:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 611) ? 241:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 612) ? 80:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 613) ? 154:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 614) ? 326:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 615) ? 394:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 616) ? 167:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 617) ? 171:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 618) ? 192:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 619) ? 275:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 620) ? 7:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 621) ? 92:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 622) ? 156:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 623) ? 339:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 624) ? 15:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 625) ? 70:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 626) ? 301:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 627) ? 314:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 628) ? 120:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 629) ? 145:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 630) ? 160:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 631) ? 337:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 632) ? 51:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 633) ? 132:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 634) ? 138:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 635) ? 227:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 636) ? 4:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 637) ? 164:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 638) ? 260:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 639) ? 291:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 640) ? 84:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 641) ? 172:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 642) ? 208:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 643) ? 233:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 644) ? 21:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 645) ? 123:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 646) ? 217:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 647) ? 303:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 648) ? 106:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 649) ? 297:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 650) ? 341:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 651) ? 397:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 652) ? 155:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 653) ? 200:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 654) ? 288:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 655) ? 363:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 656) ? 29:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 657) ? 211:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 658) ? 262:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 659) ? 378:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 660) ? 54:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 661) ? 128:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 662) ? 133:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 663) ? 269:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 664) ? 6:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 665) ? 68:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 666) ? 220:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 667) ? 362:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 668) ? 39:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 669) ? 279:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 670) ? 358:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 671) ? 367:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 672) ? 55:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 673) ? 104:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 674) ? 115:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 675) ? 263:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 676) ? 24:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 677) ? 165:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 678) ? 203:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 679) ? 302:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 680) ? 94:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 681) ? 348:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 682) ? 393:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 683) ? 395:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 684) ? 117:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 685) ? 175:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 686) ? 322:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 687) ? 381:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 688) ? 27:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 689) ? 31:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 690) ? 255:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 691) ? 366:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 692) ? 124:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 693) ? 163:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 694) ? 268:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 695) ? 390:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 696) ? 42:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 697) ? 179:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 698) ? 287:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 699) ? 321:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 700) ? 71:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 701) ? 109:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 702) ? 157:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 703) ? 284:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 704) ? 28:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 705) ? 169:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 706) ? 225:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 707) ? 232:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 708) ? 81:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 709) ? 149:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 710) ? 289:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 711) ? 374:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 712) ? 41:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 713) ? 121:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 714) ? 230:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 715) ? 305:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 716) ? 33:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 717) ? 91:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 718) ? 114:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 719) ? 216:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 720) ? 134:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 721) ? 139:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 722) ? 333:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 723) ? 357:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 724) ? 26:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 725) ? 47:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 726) ? 177:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 727) ? 259:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 728) ? 60:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 729) ? 103:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 730) ? 318:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 731) ? 338:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 732) ? 2:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 733) ? 141:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 734) ? 253:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 735) ? 282:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 736) ? 93:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 737) ? 222:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 738) ? 313:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 739) ? 316:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 740) ? 17:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 741) ? 176:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 742) ? 245:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 743) ? 370:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 744) ? 87:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 745) ? 100:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 746) ? 240:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 747) ? 265:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 748) ? 63:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 749) ? 77:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 750) ? 281:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 751) ? 349:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 752) ? 58:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 753) ? 66:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 754) ? 148:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 755) ? 306:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 756) ? 97:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 757) ? 308:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 758) ? 342:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 759) ? 355:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 760) ? 159:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 761) ? 191:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 762) ? 336:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 763) ? 345:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 764) ? 44:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 765) ? 73:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 766) ? 215:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 767) ? 309:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 768) ? 56:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 769) ? 75:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 770) ? 235:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 771) ? 307:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 772) ? 1:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 773) ? 23:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 774) ? 264:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 775) ? 386:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 776) ? 20:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 777) ? 90:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 778) ? 147:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 779) ? 237:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 780) ? 111:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 781) ? 186:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 782) ? 351:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 783) ? 369:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 784) ? 0:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 785) ? 185:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 786) ? 247:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 787) ? 340:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 788) ? 12:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 789) ? 304:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 790) ? 361:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 791) ? 380:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 792) ? 9:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 793) ? 193:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 794) ? 204:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 795) ? 311:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 796) ? 83:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 797) ? 85:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 798) ? 181:
			 /**/
			 (r_state == zStateBetaInit) & (r_counter == 799) ? 256:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1) ? 125:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 3) ? 201:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 5) ? 202:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 7) ? 203:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 9) ? 204:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 11) ? 205:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 13) ? 206:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 15) ? 207:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 17) ? 208:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 19) ? 209:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 21) ? 210:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 23) ? 211:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 25) ? 212:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 27) ? 213:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 29) ? 214:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 31) ? 215:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 33) ? 216:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 35) ? 217:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 37) ? 218:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 39) ? 219:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 41) ? 220:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 43) ? 221:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 45) ? 222:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 47) ? 223:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 49) ? 224:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 51) ? 225:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 53) ? 226:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 55) ? 227:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 57) ? 228:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 59) ? 229:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 61) ? 230:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 63) ? 231:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 65) ? 232:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 67) ? 233:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 69) ? 234:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 71) ? 235:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 73) ? 236:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 75) ? 237:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 77) ? 238:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 79) ? 239:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 81) ? 240:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 83) ? 241:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 85) ? 242:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 87) ? 243:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 89) ? 244:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 91) ? 245:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 93) ? 246:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 95) ? 247:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 97) ? 9:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 99) ? 248:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 101) ? 249:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 103) ? 250:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 105) ? 251:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 107) ? 252:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 109) ? 253:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 111) ? 254:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 113) ? 255:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 115) ? 256:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 117) ? 257:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 119) ? 258:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 121) ? 259:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 123) ? 260:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 125) ? 261:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 127) ? 262:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 129) ? 61:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 131) ? 263:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 133) ? 264:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 135) ? 265:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 137) ? 266:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 139) ? 267:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 141) ? 268:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 143) ? 269:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 145) ? 29:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 147) ? 270:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 149) ? 271:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 151) ? 272:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 153) ? 273:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 155) ? 274:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 157) ? 275:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 159) ? 276:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 161) ? 277:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 163) ? 278:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 165) ? 279:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 167) ? 280:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 169) ? 101:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 171) ? 281:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 173) ? 282:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 175) ? 283:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 177) ? 13:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 179) ? 284:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 181) ? 285:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 183) ? 286:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 185) ? 287:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 187) ? 288:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 189) ? 289:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 191) ? 290:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 193) ? 53:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 195) ? 54:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 197) ? 291:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 199) ? 292:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 201) ? 157:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 203) ? 293:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 205) ? 294:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 207) ? 295:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 209) ? 296:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 211) ? 297:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 213) ? 298:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 215) ? 299:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 217) ? 65:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 219) ? 300:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 221) ? 301:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 223) ? 302:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 225) ? 5:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 227) ? 173:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 229) ? 303:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 231) ? 304:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 233) ? 17:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 235) ? 21:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 237) ? 305:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 239) ? 306:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 241) ? 33:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 243) ? 41:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 245) ? 49:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 247) ? 307:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 249) ? 57:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 251) ? 308:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 253) ? 309:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 255) ? 310:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 257) ? 69:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 259) ? 85:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 261) ? 97:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 263) ? 311:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 265) ? 105:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 267) ? 110:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 269) ? 121:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 271) ? 312:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 273) ? 129:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 275) ? 133:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 277) ? 141:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 279) ? 313:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 281) ? 1:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 283) ? 189:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 285) ? 314:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 287) ? 315:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 289) ? 16:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 291) ? 316:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 293) ? 317:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 295) ? 318:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 297) ? 23:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 299) ? 25:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 301) ? 319:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 303) ? 320:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 305) ? 30:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 307) ? 37:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 309) ? 321:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 311) ? 322:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 313) ? 45:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 315) ? 323:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 317) ? 324:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 319) ? 325:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 321) ? 326:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 323) ? 327:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 325) ? 328:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 327) ? 329:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 329) ? 73:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 331) ? 77:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 333) ? 81:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 335) ? 330:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 337) ? 89:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 339) ? 91:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 341) ? 93:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 343) ? 331:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 345) ? 109:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 347) ? 332:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 349) ? 333:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 351) ? 334:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 353) ? 113:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 355) ? 117:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 357) ? 335:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 359) ? 336:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 361) ? 137:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 363) ? 337:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 365) ? 338:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 367) ? 339:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 369) ? 145:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 371) ? 149:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 373) ? 153:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 375) ? 340:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 377) ? 161:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 379) ? 165:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 381) ? 169:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 383) ? 341:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 385) ? 177:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 387) ? 181:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 389) ? 185:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 391) ? 342:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 393) ? 0:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 395) ? 193:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 397) ? 197:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 399) ? 343:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 401) ? 2:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 403) ? 3:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 405) ? 4:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 407) ? 344:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 409) ? 6:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 411) ? 7:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 413) ? 8:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 415) ? 345:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 417) ? 10:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 419) ? 11:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 421) ? 12:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 423) ? 346:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 425) ? 14:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 427) ? 15:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 429) ? 347:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 431) ? 348:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 433) ? 18:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 435) ? 19:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 437) ? 20:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 439) ? 349:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 441) ? 22:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 443) ? 24:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 445) ? 350:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 447) ? 351:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 449) ? 26:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 451) ? 27:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 453) ? 28:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 455) ? 352:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 457) ? 31:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 459) ? 32:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 461) ? 353:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 463) ? 354:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 465) ? 34:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 467) ? 35:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 469) ? 36:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 471) ? 355:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 473) ? 38:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 475) ? 39:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 477) ? 40:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 479) ? 356:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 481) ? 42:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 483) ? 43:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 485) ? 44:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 487) ? 357:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 489) ? 46:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 491) ? 47:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 493) ? 48:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 495) ? 358:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 497) ? 50:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 499) ? 51:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 501) ? 52:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 503) ? 359:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 505) ? 55:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 507) ? 56:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 509) ? 360:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 511) ? 361:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 513) ? 58:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 515) ? 59:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 517) ? 60:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 519) ? 362:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 521) ? 62:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 523) ? 63:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 525) ? 64:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 527) ? 363:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 529) ? 66:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 531) ? 67:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 533) ? 68:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 535) ? 364:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 537) ? 70:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 539) ? 71:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 541) ? 72:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 543) ? 365:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 545) ? 74:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 547) ? 75:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 549) ? 76:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 551) ? 366:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 553) ? 78:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 555) ? 79:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 557) ? 80:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 559) ? 367:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 561) ? 82:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 563) ? 83:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 565) ? 84:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 567) ? 368:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 569) ? 86:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 571) ? 87:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 573) ? 88:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 575) ? 369:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 577) ? 90:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 579) ? 92:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 581) ? 370:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 583) ? 371:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 585) ? 94:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 587) ? 95:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 589) ? 96:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 591) ? 372:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 593) ? 98:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 595) ? 99:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 597) ? 100:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 599) ? 373:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 601) ? 102:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 603) ? 103:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 605) ? 104:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 607) ? 374:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 609) ? 106:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 611) ? 107:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 613) ? 108:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 615) ? 375:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 617) ? 111:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 619) ? 112:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 621) ? 376:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 623) ? 377:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 625) ? 114:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 627) ? 115:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 629) ? 116:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 631) ? 378:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 633) ? 118:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 635) ? 119:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 637) ? 120:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 639) ? 379:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 641) ? 122:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 643) ? 123:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 645) ? 124:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 647) ? 380:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 649) ? 126:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 651) ? 127:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 653) ? 128:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 655) ? 381:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 657) ? 130:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 659) ? 131:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 661) ? 132:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 663) ? 382:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 665) ? 134:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 667) ? 135:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 669) ? 136:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 671) ? 383:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 673) ? 138:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 675) ? 139:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 677) ? 140:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 679) ? 384:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 681) ? 142:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 683) ? 143:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 685) ? 144:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 687) ? 385:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 689) ? 146:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 691) ? 147:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 693) ? 148:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 695) ? 386:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 697) ? 150:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 699) ? 151:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 701) ? 152:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 703) ? 387:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 705) ? 154:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 707) ? 155:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 709) ? 156:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 711) ? 388:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 713) ? 158:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 715) ? 159:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 717) ? 160:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 719) ? 389:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 721) ? 162:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 723) ? 163:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 725) ? 164:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 727) ? 390:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 729) ? 166:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 731) ? 167:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 733) ? 168:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 735) ? 391:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 737) ? 170:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 739) ? 171:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 741) ? 172:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 743) ? 392:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 745) ? 174:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 747) ? 175:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 749) ? 176:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 751) ? 393:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 753) ? 178:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 755) ? 179:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 757) ? 180:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 759) ? 394:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 761) ? 182:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 763) ? 183:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 765) ? 184:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 767) ? 395:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 769) ? 186:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 771) ? 187:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 773) ? 188:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 775) ? 396:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 777) ? 190:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 779) ? 191:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 781) ? 192:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 783) ? 397:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 785) ? 194:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 787) ? 195:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 789) ? 196:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 791) ? 398:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 793) ? 198:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 795) ? 199:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 797) ? 200:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 799) ? 399:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 801) ? 74:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 803) ? 135:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 805) ? 178:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 807) ? 325:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 809) ? 205:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 811) ? 236:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 813) ? 285:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 815) ? 335:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 817) ? 22:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 819) ? 82:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 821) ? 334:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 823) ? 391:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 825) ? 113:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 827) ? 126:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 829) ? 298:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 831) ? 329:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 833) ? 8:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 835) ? 69:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 837) ? 295:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 839) ? 385:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 841) ? 11:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 843) ? 198:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 845) ? 207:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 847) ? 332:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 849) ? 189:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 851) ? 258:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 853) ? 271:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 855) ? 346:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 857) ? 46:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 859) ? 65:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 861) ? 300:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 863) ? 347:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 865) ? 52:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 867) ? 101:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 869) ? 210:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 871) ? 376:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 873) ? 37:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 875) ? 110:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 877) ? 196:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 879) ? 257:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 881) ? 161:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 883) ? 277:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 885) ? 312:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 887) ? 356:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 889) ? 98:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 891) ? 112:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 893) ? 174:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 895) ? 317:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 897) ? 61:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 899) ? 88:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 901) ? 130:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 903) ? 250:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 905) ? 131:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 907) ? 199:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 909) ? 377:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 911) ? 399:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 913) ? 64:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 915) ? 102:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 917) ? 324:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 919) ? 368:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 921) ? 254:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 923) ? 343:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 925) ? 359:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 927) ? 372:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 929) ? 10:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 931) ? 30:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 933) ? 180:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 935) ? 243:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 937) ? 105:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 939) ? 228:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 941) ? 331:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 943) ? 365:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 945) ? 18:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 947) ? 79:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 949) ? 226:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 951) ? 296:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 953) ? 13:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 955) ? 150:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 957) ? 194:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 959) ? 280:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 961) ? 96:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 963) ? 136:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 965) ? 195:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 967) ? 315:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 969) ? 119:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 971) ? 129:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 973) ? 252:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 975) ? 353:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 977) ? 173:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 979) ? 202:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 981) ? 223:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 983) ? 389:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 985) ? 50:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 987) ? 137:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 989) ? 229:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 991) ? 272:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 993) ? 16:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 995) ? 40:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 997) ? 86:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 999) ? 293:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1001) ? 99:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1003) ? 221:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1005) ? 244:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1007) ? 267:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1009) ? 38:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1011) ? 95:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1013) ? 184:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1015) ? 327:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1017) ? 53:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1019) ? 206:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1021) ? 242:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1023) ? 248:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1025) ? 3:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1027) ? 72:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1029) ? 238:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1031) ? 383:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1033) ? 45:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1035) ? 212:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1037) ? 251:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1039) ? 379:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1041) ? 168:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1043) ? 182:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1045) ? 299:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1047) ? 392:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1049) ? 78:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1051) ? 190:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1053) ? 286:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1055) ? 384:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1057) ? 59:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1059) ? 67:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1061) ? 187:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1063) ? 354:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1065) ? 89:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1067) ? 108:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1069) ? 274:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1071) ? 375:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1073) ? 153:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1075) ? 213:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1077) ? 246:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1079) ? 398:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1081) ? 36:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1083) ? 261:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1085) ? 270:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1087) ? 283:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1089) ? 118:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1091) ? 144:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1093) ? 151:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1095) ? 371:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1097) ? 76:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1099) ? 107:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1101) ? 292:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1103) ? 330:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1105) ? 25:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1107) ? 35:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1109) ? 214:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1111) ? 294:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1113) ? 49:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1115) ? 162:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1117) ? 224:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1119) ? 382:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1121) ? 5:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1123) ? 209:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1125) ? 273:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1127) ? 344:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1129) ? 34:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1131) ? 125:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1133) ? 201:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1135) ? 319:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1137) ? 140:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1139) ? 146:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1141) ? 320:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1143) ? 388:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1145) ? 19:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1147) ? 183:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1149) ? 310:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1151) ? 373:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1153) ? 48:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1155) ? 57:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1157) ? 170:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1159) ? 234:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1161) ? 116:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1163) ? 239:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1165) ? 350:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1167) ? 364:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1169) ? 32:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1171) ? 127:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1173) ? 152:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1175) ? 328:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1177) ? 142:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1179) ? 188:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1181) ? 360:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1183) ? 396:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1185) ? 158:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1187) ? 218:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1189) ? 266:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1191) ? 352:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1193) ? 166:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1195) ? 249:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1197) ? 276:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1199) ? 323:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1201) ? 43:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1203) ? 197:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1205) ? 219:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1207) ? 290:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1209) ? 14:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1211) ? 231:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1213) ? 278:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1215) ? 387:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1217) ? 62:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1219) ? 122:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1221) ? 143:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1223) ? 241:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1225) ? 80:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1227) ? 154:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1229) ? 326:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1231) ? 394:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1233) ? 167:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1235) ? 171:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1237) ? 192:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1239) ? 275:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1241) ? 7:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1243) ? 92:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1245) ? 156:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1247) ? 339:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1249) ? 15:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1251) ? 70:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1253) ? 301:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1255) ? 314:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1257) ? 120:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1259) ? 145:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1261) ? 160:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1263) ? 337:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1265) ? 51:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1267) ? 132:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1269) ? 138:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1271) ? 227:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1273) ? 4:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1275) ? 164:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1277) ? 260:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1279) ? 291:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1281) ? 84:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1283) ? 172:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1285) ? 208:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1287) ? 233:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1289) ? 21:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1291) ? 123:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1293) ? 217:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1295) ? 303:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1297) ? 106:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1299) ? 297:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1301) ? 341:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1303) ? 397:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1305) ? 155:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1307) ? 200:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1309) ? 288:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1311) ? 363:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1313) ? 29:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1315) ? 211:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1317) ? 262:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1319) ? 378:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1321) ? 54:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1323) ? 128:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1325) ? 133:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1327) ? 269:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1329) ? 6:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1331) ? 68:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1333) ? 220:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1335) ? 362:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1337) ? 39:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1339) ? 279:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1341) ? 358:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1343) ? 367:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1345) ? 55:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1347) ? 104:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1349) ? 115:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1351) ? 263:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1353) ? 24:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1355) ? 165:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1357) ? 203:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1359) ? 302:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1361) ? 94:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1363) ? 348:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1365) ? 393:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1367) ? 395:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1369) ? 117:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1371) ? 175:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1373) ? 322:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1375) ? 381:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1377) ? 27:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1379) ? 31:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1381) ? 255:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1383) ? 366:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1385) ? 124:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1387) ? 163:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1389) ? 268:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1391) ? 390:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1393) ? 42:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1395) ? 179:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1397) ? 287:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1399) ? 321:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1401) ? 71:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1403) ? 109:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1405) ? 157:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1407) ? 284:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1409) ? 28:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1411) ? 169:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1413) ? 225:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1415) ? 232:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1417) ? 81:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1419) ? 149:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1421) ? 289:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1423) ? 374:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1425) ? 41:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1427) ? 121:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1429) ? 230:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1431) ? 305:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1433) ? 33:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1435) ? 91:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1437) ? 114:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1439) ? 216:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1441) ? 134:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1443) ? 139:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1445) ? 333:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1447) ? 357:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1449) ? 26:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1451) ? 47:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1453) ? 177:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1455) ? 259:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1457) ? 60:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1459) ? 103:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1461) ? 318:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1463) ? 338:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1465) ? 2:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1467) ? 141:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1469) ? 253:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1471) ? 282:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1473) ? 93:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1475) ? 222:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1477) ? 313:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1479) ? 316:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1481) ? 17:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1483) ? 176:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1485) ? 245:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1487) ? 370:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1489) ? 87:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1491) ? 100:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1493) ? 240:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1495) ? 265:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1497) ? 63:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1499) ? 77:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1501) ? 281:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1503) ? 349:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1505) ? 58:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1507) ? 66:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1509) ? 148:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1511) ? 306:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1513) ? 97:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1515) ? 308:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1517) ? 342:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1519) ? 355:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1521) ? 159:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1523) ? 191:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1525) ? 336:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1527) ? 345:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1529) ? 44:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1531) ? 73:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1533) ? 215:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1535) ? 309:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1537) ? 56:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1539) ? 75:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1541) ? 235:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1543) ? 307:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1545) ? 1:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1547) ? 23:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1549) ? 264:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1551) ? 386:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1553) ? 20:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1555) ? 90:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1557) ? 147:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1559) ? 237:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1561) ? 111:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1563) ? 186:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1565) ? 351:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1567) ? 369:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1569) ? 0:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1571) ? 185:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1573) ? 247:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1575) ? 340:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1577) ? 12:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1579) ? 304:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1581) ? 361:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1583) ? 380:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1585) ? 9:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1587) ? 193:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1589) ? 204:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1591) ? 311:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1593) ? 83:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1595) ? 85:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1597) ? 181:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/ 
			 (r_state == zStateColumn) & (r_counter == 1599) ? 256:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 2 & r_state==zStateEstimate) ? 0:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 5 & r_state==zStateEstimate) ? 1:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 8 & r_state==zStateEstimate) ? 2:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 11 & r_state==zStateEstimate) ? 3:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 14 & r_state==zStateEstimate) ? 4:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 17 & r_state==zStateEstimate) ? 5:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 20 & r_state==zStateEstimate) ? 6:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 23 & r_state==zStateEstimate) ? 7:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 26 & r_state==zStateEstimate) ? 8:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 29 & r_state==zStateEstimate) ? 9:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 32 & r_state==zStateEstimate) ? 10:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 35 & r_state==zStateEstimate) ? 11:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 38 & r_state==zStateEstimate) ? 12:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 41 & r_state==zStateEstimate) ? 13:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 44 & r_state==zStateEstimate) ? 14:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 47 & r_state==zStateEstimate) ? 15:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 50 & r_state==zStateEstimate) ? 16:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 53 & r_state==zStateEstimate) ? 17:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 56 & r_state==zStateEstimate) ? 18:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 59 & r_state==zStateEstimate) ? 19:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 62 & r_state==zStateEstimate) ? 20:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 65 & r_state==zStateEstimate) ? 21:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 68 & r_state==zStateEstimate) ? 22:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 71 & r_state==zStateEstimate) ? 23:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 74 & r_state==zStateEstimate) ? 24:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 77 & r_state==zStateEstimate) ? 25:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 80 & r_state==zStateEstimate) ? 26:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 83 & r_state==zStateEstimate) ? 27:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 86 & r_state==zStateEstimate) ? 28:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 89 & r_state==zStateEstimate) ? 29:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 92 & r_state==zStateEstimate) ? 30:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 95 & r_state==zStateEstimate) ? 31:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 98 & r_state==zStateEstimate) ? 32:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 101 & r_state==zStateEstimate) ? 33:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 104 & r_state==zStateEstimate) ? 34:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 107 & r_state==zStateEstimate) ? 35:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 110 & r_state==zStateEstimate) ? 36:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 113 & r_state==zStateEstimate) ? 37:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 116 & r_state==zStateEstimate) ? 38:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 119 & r_state==zStateEstimate) ? 39:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 122 & r_state==zStateEstimate) ? 40:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 125 & r_state==zStateEstimate) ? 41:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 128 & r_state==zStateEstimate) ? 42:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 131 & r_state==zStateEstimate) ? 43:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 134 & r_state==zStateEstimate) ? 44:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 137 & r_state==zStateEstimate) ? 45:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 140 & r_state==zStateEstimate) ? 46:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 143 & r_state==zStateEstimate) ? 47:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 146 & r_state==zStateEstimate) ? 48:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 149 & r_state==zStateEstimate) ? 49:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 152 & r_state==zStateEstimate) ? 50:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 155 & r_state==zStateEstimate) ? 51:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 158 & r_state==zStateEstimate) ? 52:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 161 & r_state==zStateEstimate) ? 53:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 164 & r_state==zStateEstimate) ? 54:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 167 & r_state==zStateEstimate) ? 55:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 170 & r_state==zStateEstimate) ? 56:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 173 & r_state==zStateEstimate) ? 57:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 176 & r_state==zStateEstimate) ? 58:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 179 & r_state==zStateEstimate) ? 59:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 182 & r_state==zStateEstimate) ? 60:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 185 & r_state==zStateEstimate) ? 61:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 188 & r_state==zStateEstimate) ? 62:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 191 & r_state==zStateEstimate) ? 63:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 194 & r_state==zStateEstimate) ? 64:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 197 & r_state==zStateEstimate) ? 65:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 200 & r_state==zStateEstimate) ? 66:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 203 & r_state==zStateEstimate) ? 67:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 206 & r_state==zStateEstimate) ? 68:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 209 & r_state==zStateEstimate) ? 69:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 212 & r_state==zStateEstimate) ? 70:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 215 & r_state==zStateEstimate) ? 71:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 218 & r_state==zStateEstimate) ? 72:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 221 & r_state==zStateEstimate) ? 73:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 224 & r_state==zStateEstimate) ? 74:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 227 & r_state==zStateEstimate) ? 75:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 230 & r_state==zStateEstimate) ? 76:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 233 & r_state==zStateEstimate) ? 77:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 236 & r_state==zStateEstimate) ? 78:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 239 & r_state==zStateEstimate) ? 79:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 242 & r_state==zStateEstimate) ? 80:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 245 & r_state==zStateEstimate) ? 81:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 248 & r_state==zStateEstimate) ? 82:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 251 & r_state==zStateEstimate) ? 83:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 254 & r_state==zStateEstimate) ? 84:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 257 & r_state==zStateEstimate) ? 85:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 260 & r_state==zStateEstimate) ? 86:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 263 & r_state==zStateEstimate) ? 87:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 266 & r_state==zStateEstimate) ? 88:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 269 & r_state==zStateEstimate) ? 89:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 272 & r_state==zStateEstimate) ? 90:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 275 & r_state==zStateEstimate) ? 91:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 278 & r_state==zStateEstimate) ? 92:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 281 & r_state==zStateEstimate) ? 93:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 284 & r_state==zStateEstimate) ? 94:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 287 & r_state==zStateEstimate) ? 95:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 290 & r_state==zStateEstimate) ? 96:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 293 & r_state==zStateEstimate) ? 97:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 296 & r_state==zStateEstimate) ? 98:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 299 & r_state==zStateEstimate) ? 99:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 302 & r_state==zStateEstimate) ? 100:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 305 & r_state==zStateEstimate) ? 101:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 308 & r_state==zStateEstimate) ? 102:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 311 & r_state==zStateEstimate) ? 103:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 314 & r_state==zStateEstimate) ? 104:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 317 & r_state==zStateEstimate) ? 105:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 320 & r_state==zStateEstimate) ? 106:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 323 & r_state==zStateEstimate) ? 107:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 326 & r_state==zStateEstimate) ? 108:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 329 & r_state==zStateEstimate) ? 109:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 332 & r_state==zStateEstimate) ? 110:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 335 & r_state==zStateEstimate) ? 111:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 338 & r_state==zStateEstimate) ? 112:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 341 & r_state==zStateEstimate) ? 113:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 344 & r_state==zStateEstimate) ? 114:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 347 & r_state==zStateEstimate) ? 115:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 350 & r_state==zStateEstimate) ? 116:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 353 & r_state==zStateEstimate) ? 117:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 356 & r_state==zStateEstimate) ? 118:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 359 & r_state==zStateEstimate) ? 119:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 362 & r_state==zStateEstimate) ? 120:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 365 & r_state==zStateEstimate) ? 121:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 368 & r_state==zStateEstimate) ? 122:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 371 & r_state==zStateEstimate) ? 123:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 374 & r_state==zStateEstimate) ? 124:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 377 & r_state==zStateEstimate) ? 125:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 380 & r_state==zStateEstimate) ? 126:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 383 & r_state==zStateEstimate) ? 127:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 386 & r_state==zStateEstimate) ? 128:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 389 & r_state==zStateEstimate) ? 129:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 392 & r_state==zStateEstimate) ? 130:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 395 & r_state==zStateEstimate) ? 131:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 398 & r_state==zStateEstimate) ? 132:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 401 & r_state==zStateEstimate) ? 133:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 404 & r_state==zStateEstimate) ? 134:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 407 & r_state==zStateEstimate) ? 135:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 410 & r_state==zStateEstimate) ? 136:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 413 & r_state==zStateEstimate) ? 137:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 416 & r_state==zStateEstimate) ? 138:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 419 & r_state==zStateEstimate) ? 139:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 422 & r_state==zStateEstimate) ? 140:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 425 & r_state==zStateEstimate) ? 141:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 428 & r_state==zStateEstimate) ? 142:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 431 & r_state==zStateEstimate) ? 143:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 434 & r_state==zStateEstimate) ? 144:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 437 & r_state==zStateEstimate) ? 145:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 440 & r_state==zStateEstimate) ? 146:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 443 & r_state==zStateEstimate) ? 147:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 446 & r_state==zStateEstimate) ? 148:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 449 & r_state==zStateEstimate) ? 149:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 452 & r_state==zStateEstimate) ? 150:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 455 & r_state==zStateEstimate) ? 151:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 458 & r_state==zStateEstimate) ? 152:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 461 & r_state==zStateEstimate) ? 153:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 464 & r_state==zStateEstimate) ? 154:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 467 & r_state==zStateEstimate) ? 155:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 470 & r_state==zStateEstimate) ? 156:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 473 & r_state==zStateEstimate) ? 157:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 476 & r_state==zStateEstimate) ? 158:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 479 & r_state==zStateEstimate) ? 159:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 482 & r_state==zStateEstimate) ? 160:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 485 & r_state==zStateEstimate) ? 161:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 488 & r_state==zStateEstimate) ? 162:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 491 & r_state==zStateEstimate) ? 163:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 494 & r_state==zStateEstimate) ? 164:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 497 & r_state==zStateEstimate) ? 165:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 500 & r_state==zStateEstimate) ? 166:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 503 & r_state==zStateEstimate) ? 167:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 506 & r_state==zStateEstimate) ? 168:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 509 & r_state==zStateEstimate) ? 169:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 512 & r_state==zStateEstimate) ? 170:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 515 & r_state==zStateEstimate) ? 171:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 518 & r_state==zStateEstimate) ? 172:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 521 & r_state==zStateEstimate) ? 173:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 524 & r_state==zStateEstimate) ? 174:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 527 & r_state==zStateEstimate) ? 175:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 530 & r_state==zStateEstimate) ? 176:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 533 & r_state==zStateEstimate) ? 177:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 536 & r_state==zStateEstimate) ? 178:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 539 & r_state==zStateEstimate) ? 179:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 542 & r_state==zStateEstimate) ? 180:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 545 & r_state==zStateEstimate) ? 181:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 548 & r_state==zStateEstimate) ? 182:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 551 & r_state==zStateEstimate) ? 183:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 554 & r_state==zStateEstimate) ? 184:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 557 & r_state==zStateEstimate) ? 185:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 560 & r_state==zStateEstimate) ? 186:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 563 & r_state==zStateEstimate) ? 187:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 566 & r_state==zStateEstimate) ? 188:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 569 & r_state==zStateEstimate) ? 189:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 572 & r_state==zStateEstimate) ? 190:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 575 & r_state==zStateEstimate) ? 191:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 578 & r_state==zStateEstimate) ? 192:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 581 & r_state==zStateEstimate) ? 193:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 584 & r_state==zStateEstimate) ? 194:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 587 & r_state==zStateEstimate) ? 195:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 590 & r_state==zStateEstimate) ? 196:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 593 & r_state==zStateEstimate) ? 197:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 596 & r_state==zStateEstimate) ? 198:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 599 & r_state==zStateEstimate) ? 199:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 602 & r_state==zStateEstimate) ? 200:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 605 & r_state==zStateEstimate) ? 201:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 608 & r_state==zStateEstimate) ? 202:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 611 & r_state==zStateEstimate) ? 203:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 614 & r_state==zStateEstimate) ? 204:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 617 & r_state==zStateEstimate) ? 205:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 620 & r_state==zStateEstimate) ? 206:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 623 & r_state==zStateEstimate) ? 207:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 626 & r_state==zStateEstimate) ? 208:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 629 & r_state==zStateEstimate) ? 209:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 632 & r_state==zStateEstimate) ? 210:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 635 & r_state==zStateEstimate) ? 211:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 638 & r_state==zStateEstimate) ? 212:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 641 & r_state==zStateEstimate) ? 213:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 644 & r_state==zStateEstimate) ? 214:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 647 & r_state==zStateEstimate) ? 215:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 650 & r_state==zStateEstimate) ? 216:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 653 & r_state==zStateEstimate) ? 217:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 656 & r_state==zStateEstimate) ? 218:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 659 & r_state==zStateEstimate) ? 219:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 662 & r_state==zStateEstimate) ? 220:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 665 & r_state==zStateEstimate) ? 221:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 668 & r_state==zStateEstimate) ? 222:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 671 & r_state==zStateEstimate) ? 223:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 674 & r_state==zStateEstimate) ? 224:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 677 & r_state==zStateEstimate) ? 225:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 680 & r_state==zStateEstimate) ? 226:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 683 & r_state==zStateEstimate) ? 227:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 686 & r_state==zStateEstimate) ? 228:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 689 & r_state==zStateEstimate) ? 229:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 692 & r_state==zStateEstimate) ? 230:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 695 & r_state==zStateEstimate) ? 231:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 698 & r_state==zStateEstimate) ? 232:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 701 & r_state==zStateEstimate) ? 233:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 704 & r_state==zStateEstimate) ? 234:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 707 & r_state==zStateEstimate) ? 235:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 710 & r_state==zStateEstimate) ? 236:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 713 & r_state==zStateEstimate) ? 237:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 716 & r_state==zStateEstimate) ? 238:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 719 & r_state==zStateEstimate) ? 239:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 722 & r_state==zStateEstimate) ? 240:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 725 & r_state==zStateEstimate) ? 241:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 728 & r_state==zStateEstimate) ? 242:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 731 & r_state==zStateEstimate) ? 243:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 734 & r_state==zStateEstimate) ? 244:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 737 & r_state==zStateEstimate) ? 245:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 740 & r_state==zStateEstimate) ? 246:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 743 & r_state==zStateEstimate) ? 247:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 746 & r_state==zStateEstimate) ? 248:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 749 & r_state==zStateEstimate) ? 249:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 752 & r_state==zStateEstimate) ? 250:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 755 & r_state==zStateEstimate) ? 251:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 758 & r_state==zStateEstimate) ? 252:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 761 & r_state==zStateEstimate) ? 253:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 764 & r_state==zStateEstimate) ? 254:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 767 & r_state==zStateEstimate) ? 255:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 770 & r_state==zStateEstimate) ? 256:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 773 & r_state==zStateEstimate) ? 257:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 776 & r_state==zStateEstimate) ? 258:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 779 & r_state==zStateEstimate) ? 259:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 782 & r_state==zStateEstimate) ? 260:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 785 & r_state==zStateEstimate) ? 261:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 788 & r_state==zStateEstimate) ? 262:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 791 & r_state==zStateEstimate) ? 263:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 794 & r_state==zStateEstimate) ? 264:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 797 & r_state==zStateEstimate) ? 265:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 800 & r_state==zStateEstimate) ? 266:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 803 & r_state==zStateEstimate) ? 267:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 806 & r_state==zStateEstimate) ? 268:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 809 & r_state==zStateEstimate) ? 269:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 812 & r_state==zStateEstimate) ? 270:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 815 & r_state==zStateEstimate) ? 271:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 818 & r_state==zStateEstimate) ? 272:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 821 & r_state==zStateEstimate) ? 273:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 824 & r_state==zStateEstimate) ? 274:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 827 & r_state==zStateEstimate) ? 275:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 830 & r_state==zStateEstimate) ? 276:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 833 & r_state==zStateEstimate) ? 277:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 836 & r_state==zStateEstimate) ? 278:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 839 & r_state==zStateEstimate) ? 279:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 842 & r_state==zStateEstimate) ? 280:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 845 & r_state==zStateEstimate) ? 281:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 848 & r_state==zStateEstimate) ? 282:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 851 & r_state==zStateEstimate) ? 283:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 854 & r_state==zStateEstimate) ? 284:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 857 & r_state==zStateEstimate) ? 285:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 860 & r_state==zStateEstimate) ? 286:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 863 & r_state==zStateEstimate) ? 287:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 866 & r_state==zStateEstimate) ? 288:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 869 & r_state==zStateEstimate) ? 289:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 872 & r_state==zStateEstimate) ? 290:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 875 & r_state==zStateEstimate) ? 291:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 878 & r_state==zStateEstimate) ? 292:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 881 & r_state==zStateEstimate) ? 293:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 884 & r_state==zStateEstimate) ? 294:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 887 & r_state==zStateEstimate) ? 295:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 890 & r_state==zStateEstimate) ? 296:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 893 & r_state==zStateEstimate) ? 297:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 896 & r_state==zStateEstimate) ? 298:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 899 & r_state==zStateEstimate) ? 299:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 902 & r_state==zStateEstimate) ? 300:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 905 & r_state==zStateEstimate) ? 301:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 908 & r_state==zStateEstimate) ? 302:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 911 & r_state==zStateEstimate) ? 303:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 914 & r_state==zStateEstimate) ? 304:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 917 & r_state==zStateEstimate) ? 305:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 920 & r_state==zStateEstimate) ? 306:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 923 & r_state==zStateEstimate) ? 307:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 926 & r_state==zStateEstimate) ? 308:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 929 & r_state==zStateEstimate) ? 309:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 932 & r_state==zStateEstimate) ? 310:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 935 & r_state==zStateEstimate) ? 311:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 938 & r_state==zStateEstimate) ? 312:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 941 & r_state==zStateEstimate) ? 313:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 944 & r_state==zStateEstimate) ? 314:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 947 & r_state==zStateEstimate) ? 315:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 950 & r_state==zStateEstimate) ? 316:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 953 & r_state==zStateEstimate) ? 317:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 956 & r_state==zStateEstimate) ? 318:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 959 & r_state==zStateEstimate) ? 319:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 962 & r_state==zStateEstimate) ? 320:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 965 & r_state==zStateEstimate) ? 321:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 968 & r_state==zStateEstimate) ? 322:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 971 & r_state==zStateEstimate) ? 323:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 974 & r_state==zStateEstimate) ? 324:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 977 & r_state==zStateEstimate) ? 325:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 980 & r_state==zStateEstimate) ? 326:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 983 & r_state==zStateEstimate) ? 327:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 986 & r_state==zStateEstimate) ? 328:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 989 & r_state==zStateEstimate) ? 329:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 992 & r_state==zStateEstimate) ? 330:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 995 & r_state==zStateEstimate) ? 331:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 998 & r_state==zStateEstimate) ? 332:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1001 & r_state==zStateEstimate) ? 333:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1004 & r_state==zStateEstimate) ? 334:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1007 & r_state==zStateEstimate) ? 335:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1010 & r_state==zStateEstimate) ? 336:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1013 & r_state==zStateEstimate) ? 337:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1016 & r_state==zStateEstimate) ? 338:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1019 & r_state==zStateEstimate) ? 339:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1022 & r_state==zStateEstimate) ? 340:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1025 & r_state==zStateEstimate) ? 341:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1028 & r_state==zStateEstimate) ? 342:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1031 & r_state==zStateEstimate) ? 343:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1034 & r_state==zStateEstimate) ? 344:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1037 & r_state==zStateEstimate) ? 345:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1040 & r_state==zStateEstimate) ? 346:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1043 & r_state==zStateEstimate) ? 347:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1046 & r_state==zStateEstimate) ? 348:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1049 & r_state==zStateEstimate) ? 349:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1052 & r_state==zStateEstimate) ? 350:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1055 & r_state==zStateEstimate) ? 351:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1058 & r_state==zStateEstimate) ? 352:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1061 & r_state==zStateEstimate) ? 353:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1064 & r_state==zStateEstimate) ? 354:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1067 & r_state==zStateEstimate) ? 355:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1070 & r_state==zStateEstimate) ? 356:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1073 & r_state==zStateEstimate) ? 357:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1076 & r_state==zStateEstimate) ? 358:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1079 & r_state==zStateEstimate) ? 359:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1082 & r_state==zStateEstimate) ? 360:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1085 & r_state==zStateEstimate) ? 361:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1088 & r_state==zStateEstimate) ? 362:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1091 & r_state==zStateEstimate) ? 363:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1094 & r_state==zStateEstimate) ? 364:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1097 & r_state==zStateEstimate) ? 365:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1100 & r_state==zStateEstimate) ? 366:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1103 & r_state==zStateEstimate) ? 367:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1106 & r_state==zStateEstimate) ? 368:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1109 & r_state==zStateEstimate) ? 369:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1112 & r_state==zStateEstimate) ? 370:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1115 & r_state==zStateEstimate) ? 371:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1118 & r_state==zStateEstimate) ? 372:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1121 & r_state==zStateEstimate) ? 373:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1124 & r_state==zStateEstimate) ? 374:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1127 & r_state==zStateEstimate) ? 375:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1130 & r_state==zStateEstimate) ? 376:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1133 & r_state==zStateEstimate) ? 377:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1136 & r_state==zStateEstimate) ? 378:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1139 & r_state==zStateEstimate) ? 379:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1142 & r_state==zStateEstimate) ? 380:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1145 & r_state==zStateEstimate) ? 381:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1148 & r_state==zStateEstimate) ? 382:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1151 & r_state==zStateEstimate) ? 383:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1154 & r_state==zStateEstimate) ? 384:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1157 & r_state==zStateEstimate) ? 385:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1160 & r_state==zStateEstimate) ? 386:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1163 & r_state==zStateEstimate) ? 387:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1166 & r_state==zStateEstimate) ? 388:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1169 & r_state==zStateEstimate) ? 389:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1172 & r_state==zStateEstimate) ? 390:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1175 & r_state==zStateEstimate) ? 391:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1178 & r_state==zStateEstimate) ? 392:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1181 & r_state==zStateEstimate) ? 393:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1184 & r_state==zStateEstimate) ? 394:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1187 & r_state==zStateEstimate) ? 395:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1190 & r_state==zStateEstimate) ? 396:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1193 & r_state==zStateEstimate) ? 397:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1196 & r_state==zStateEstimate) ? 398:
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 /**/
			 (r_counter == 1199 & r_state==zStateEstimate) ? 399:
			 /**/
			 /**/
			 0;
   assign i_wdata_lambda=/**/
		  (r_counter==0) ? i_data[15:0]:
		  /**/
		  (r_counter==1) ? i_data[15:0]:
		  /**/
		  (r_counter==2) ? i_data[15:0]:
		  /**/
		  (r_counter==3) ? i_data[15:0]:
		  /**/
		  (r_counter==4) ? i_data[15:0]:
		  /**/
		  (r_counter==5) ? i_data[15:0]:
		  /**/
		  (r_counter==6) ? i_data[15:0]:
		  /**/
		  (r_counter==7) ? i_data[15:0]:
		  /**/
		  (r_counter==8) ? i_data[15:0]:
		  /**/
		  (r_counter==9) ? i_data[15:0]:
		  /**/
		  (r_counter==10) ? i_data[15:0]:
		  /**/
		  (r_counter==11) ? i_data[15:0]:
		  /**/
		  (r_counter==12) ? i_data[15:0]:
		  /**/
		  (r_counter==13) ? i_data[15:0]:
		  /**/
		  (r_counter==14) ? i_data[15:0]:
		  /**/
		  (r_counter==15) ? i_data[15:0]:
		  /**/
		  (r_counter==16) ? i_data[15:0]:
		  /**/
		  (r_counter==17) ? i_data[15:0]:
		  /**/
		  (r_counter==18) ? i_data[15:0]:
		  /**/
		  (r_counter==19) ? i_data[15:0]:
		  /**/
		  (r_counter==20) ? i_data[15:0]:
		  /**/
		  (r_counter==21) ? i_data[15:0]:
		  /**/
		  (r_counter==22) ? i_data[15:0]:
		  /**/
		  (r_counter==23) ? i_data[15:0]:
		  /**/
		  (r_counter==24) ? i_data[15:0]:
		  /**/
		  (r_counter==25) ? i_data[15:0]:
		  /**/
		  (r_counter==26) ? i_data[15:0]:
		  /**/
		  (r_counter==27) ? i_data[15:0]:
		  /**/
		  (r_counter==28) ? i_data[15:0]:
		  /**/
		  (r_counter==29) ? i_data[15:0]:
		  /**/
		  (r_counter==30) ? i_data[15:0]:
		  /**/
		  (r_counter==31) ? i_data[15:0]:
		  /**/
		  (r_counter==32) ? i_data[15:0]:
		  /**/
		  (r_counter==33) ? i_data[15:0]:
		  /**/
		  (r_counter==34) ? i_data[15:0]:
		  /**/
		  (r_counter==35) ? i_data[15:0]:
		  /**/
		  (r_counter==36) ? i_data[15:0]:
		  /**/
		  (r_counter==37) ? i_data[15:0]:
		  /**/
		  (r_counter==38) ? i_data[15:0]:
		  /**/
		  (r_counter==39) ? i_data[15:0]:
		  /**/
		  (r_counter==40) ? i_data[15:0]:
		  /**/
		  (r_counter==41) ? i_data[15:0]:
		  /**/
		  (r_counter==42) ? i_data[15:0]:
		  /**/
		  (r_counter==43) ? i_data[15:0]:
		  /**/
		  (r_counter==44) ? i_data[15:0]:
		  /**/
		  (r_counter==45) ? i_data[15:0]:
		  /**/
		  (r_counter==46) ? i_data[15:0]:
		  /**/
		  (r_counter==47) ? i_data[15:0]:
		  /**/
		  (r_counter==48) ? i_data[15:0]:
		  /**/
		  (r_counter==49) ? i_data[15:0]:
		  /**/
		  (r_counter==50) ? i_data[15:0]:
		  /**/
		  (r_counter==51) ? i_data[15:0]:
		  /**/
		  (r_counter==52) ? i_data[15:0]:
		  /**/
		  (r_counter==53) ? i_data[15:0]:
		  /**/
		  (r_counter==54) ? i_data[15:0]:
		  /**/
		  (r_counter==55) ? i_data[15:0]:
		  /**/
		  (r_counter==56) ? i_data[15:0]:
		  /**/
		  (r_counter==57) ? i_data[15:0]:
		  /**/
		  (r_counter==58) ? i_data[15:0]:
		  /**/
		  (r_counter==59) ? i_data[15:0]:
		  /**/
		  (r_counter==60) ? i_data[15:0]:
		  /**/
		  (r_counter==61) ? i_data[15:0]:
		  /**/
		  (r_counter==62) ? i_data[15:0]:
		  /**/
		  (r_counter==63) ? i_data[15:0]:
		  /**/
		  (r_counter==64) ? i_data[15:0]:
		  /**/
		  (r_counter==65) ? i_data[15:0]:
		  /**/
		  (r_counter==66) ? i_data[15:0]:
		  /**/
		  (r_counter==67) ? i_data[15:0]:
		  /**/
		  (r_counter==68) ? i_data[15:0]:
		  /**/
		  (r_counter==69) ? i_data[15:0]:
		  /**/
		  (r_counter==70) ? i_data[15:0]:
		  /**/
		  (r_counter==71) ? i_data[15:0]:
		  /**/
		  (r_counter==72) ? i_data[15:0]:
		  /**/
		  (r_counter==73) ? i_data[15:0]:
		  /**/
		  (r_counter==74) ? i_data[15:0]:
		  /**/
		  (r_counter==75) ? i_data[15:0]:
		  /**/
		  (r_counter==76) ? i_data[15:0]:
		  /**/
		  (r_counter==77) ? i_data[15:0]:
		  /**/
		  (r_counter==78) ? i_data[15:0]:
		  /**/
		  (r_counter==79) ? i_data[15:0]:
		  /**/
		  (r_counter==80) ? i_data[15:0]:
		  /**/
		  (r_counter==81) ? i_data[15:0]:
		  /**/
		  (r_counter==82) ? i_data[15:0]:
		  /**/
		  (r_counter==83) ? i_data[15:0]:
		  /**/
		  (r_counter==84) ? i_data[15:0]:
		  /**/
		  (r_counter==85) ? i_data[15:0]:
		  /**/
		  (r_counter==86) ? i_data[15:0]:
		  /**/
		  (r_counter==87) ? i_data[15:0]:
		  /**/
		  (r_counter==88) ? i_data[15:0]:
		  /**/
		  (r_counter==89) ? i_data[15:0]:
		  /**/
		  (r_counter==90) ? i_data[15:0]:
		  /**/
		  (r_counter==91) ? i_data[15:0]:
		  /**/
		  (r_counter==92) ? i_data[15:0]:
		  /**/
		  (r_counter==93) ? i_data[15:0]:
		  /**/
		  (r_counter==94) ? i_data[15:0]:
		  /**/
		  (r_counter==95) ? i_data[15:0]:
		  /**/
		  (r_counter==96) ? i_data[15:0]:
		  /**/
		  (r_counter==97) ? i_data[15:0]:
		  /**/
		  (r_counter==98) ? i_data[15:0]:
		  /**/
		  (r_counter==99) ? i_data[15:0]:
		  /**/
		  (r_counter==100) ? i_data[15:0]:
		  /**/
		  (r_counter==101) ? i_data[15:0]:
		  /**/
		  (r_counter==102) ? i_data[15:0]:
		  /**/
		  (r_counter==103) ? i_data[15:0]:
		  /**/
		  (r_counter==104) ? i_data[15:0]:
		  /**/
		  (r_counter==105) ? i_data[15:0]:
		  /**/
		  (r_counter==106) ? i_data[15:0]:
		  /**/
		  (r_counter==107) ? i_data[15:0]:
		  /**/
		  (r_counter==108) ? i_data[15:0]:
		  /**/
		  (r_counter==109) ? i_data[15:0]:
		  /**/
		  (r_counter==110) ? i_data[15:0]:
		  /**/
		  (r_counter==111) ? i_data[15:0]:
		  /**/
		  (r_counter==112) ? i_data[15:0]:
		  /**/
		  (r_counter==113) ? i_data[15:0]:
		  /**/
		  (r_counter==114) ? i_data[15:0]:
		  /**/
		  (r_counter==115) ? i_data[15:0]:
		  /**/
		  (r_counter==116) ? i_data[15:0]:
		  /**/
		  (r_counter==117) ? i_data[15:0]:
		  /**/
		  (r_counter==118) ? i_data[15:0]:
		  /**/
		  (r_counter==119) ? i_data[15:0]:
		  /**/
		  (r_counter==120) ? i_data[15:0]:
		  /**/
		  (r_counter==121) ? i_data[15:0]:
		  /**/
		  (r_counter==122) ? i_data[15:0]:
		  /**/
		  (r_counter==123) ? i_data[15:0]:
		  /**/
		  (r_counter==124) ? i_data[15:0]:
		  /**/
		  (r_counter==125) ? i_data[15:0]:
		  /**/
		  (r_counter==126) ? i_data[15:0]:
		  /**/
		  (r_counter==127) ? i_data[15:0]:
		  /**/
		  (r_counter==128) ? i_data[15:0]:
		  /**/
		  (r_counter==129) ? i_data[15:0]:
		  /**/
		  (r_counter==130) ? i_data[15:0]:
		  /**/
		  (r_counter==131) ? i_data[15:0]:
		  /**/
		  (r_counter==132) ? i_data[15:0]:
		  /**/
		  (r_counter==133) ? i_data[15:0]:
		  /**/
		  (r_counter==134) ? i_data[15:0]:
		  /**/
		  (r_counter==135) ? i_data[15:0]:
		  /**/
		  (r_counter==136) ? i_data[15:0]:
		  /**/
		  (r_counter==137) ? i_data[15:0]:
		  /**/
		  (r_counter==138) ? i_data[15:0]:
		  /**/
		  (r_counter==139) ? i_data[15:0]:
		  /**/
		  (r_counter==140) ? i_data[15:0]:
		  /**/
		  (r_counter==141) ? i_data[15:0]:
		  /**/
		  (r_counter==142) ? i_data[15:0]:
		  /**/
		  (r_counter==143) ? i_data[15:0]:
		  /**/
		  (r_counter==144) ? i_data[15:0]:
		  /**/
		  (r_counter==145) ? i_data[15:0]:
		  /**/
		  (r_counter==146) ? i_data[15:0]:
		  /**/
		  (r_counter==147) ? i_data[15:0]:
		  /**/
		  (r_counter==148) ? i_data[15:0]:
		  /**/
		  (r_counter==149) ? i_data[15:0]:
		  /**/
		  (r_counter==150) ? i_data[15:0]:
		  /**/
		  (r_counter==151) ? i_data[15:0]:
		  /**/
		  (r_counter==152) ? i_data[15:0]:
		  /**/
		  (r_counter==153) ? i_data[15:0]:
		  /**/
		  (r_counter==154) ? i_data[15:0]:
		  /**/
		  (r_counter==155) ? i_data[15:0]:
		  /**/
		  (r_counter==156) ? i_data[15:0]:
		  /**/
		  (r_counter==157) ? i_data[15:0]:
		  /**/
		  (r_counter==158) ? i_data[15:0]:
		  /**/
		  (r_counter==159) ? i_data[15:0]:
		  /**/
		  (r_counter==160) ? i_data[15:0]:
		  /**/
		  (r_counter==161) ? i_data[15:0]:
		  /**/
		  (r_counter==162) ? i_data[15:0]:
		  /**/
		  (r_counter==163) ? i_data[15:0]:
		  /**/
		  (r_counter==164) ? i_data[15:0]:
		  /**/
		  (r_counter==165) ? i_data[15:0]:
		  /**/
		  (r_counter==166) ? i_data[15:0]:
		  /**/
		  (r_counter==167) ? i_data[15:0]:
		  /**/
		  (r_counter==168) ? i_data[15:0]:
		  /**/
		  (r_counter==169) ? i_data[15:0]:
		  /**/
		  (r_counter==170) ? i_data[15:0]:
		  /**/
		  (r_counter==171) ? i_data[15:0]:
		  /**/
		  (r_counter==172) ? i_data[15:0]:
		  /**/
		  (r_counter==173) ? i_data[15:0]:
		  /**/
		  (r_counter==174) ? i_data[15:0]:
		  /**/
		  (r_counter==175) ? i_data[15:0]:
		  /**/
		  (r_counter==176) ? i_data[15:0]:
		  /**/
		  (r_counter==177) ? i_data[15:0]:
		  /**/
		  (r_counter==178) ? i_data[15:0]:
		  /**/
		  (r_counter==179) ? i_data[15:0]:
		  /**/
		  (r_counter==180) ? i_data[15:0]:
		  /**/
		  (r_counter==181) ? i_data[15:0]:
		  /**/
		  (r_counter==182) ? i_data[15:0]:
		  /**/
		  (r_counter==183) ? i_data[15:0]:
		  /**/
		  (r_counter==184) ? i_data[15:0]:
		  /**/
		  (r_counter==185) ? i_data[15:0]:
		  /**/
		  (r_counter==186) ? i_data[15:0]:
		  /**/
		  (r_counter==187) ? i_data[15:0]:
		  /**/
		  (r_counter==188) ? i_data[15:0]:
		  /**/
		  (r_counter==189) ? i_data[15:0]:
		  /**/
		  (r_counter==190) ? i_data[15:0]:
		  /**/
		  (r_counter==191) ? i_data[15:0]:
		  /**/
		  (r_counter==192) ? i_data[15:0]:
		  /**/
		  (r_counter==193) ? i_data[15:0]:
		  /**/
		  (r_counter==194) ? i_data[15:0]:
		  /**/
		  (r_counter==195) ? i_data[15:0]:
		  /**/
		  (r_counter==196) ? i_data[15:0]:
		  /**/
		  (r_counter==197) ? i_data[15:0]:
		  /**/
		  (r_counter==198) ? i_data[15:0]:
		  /**/
		  (r_counter==199) ? i_data[15:0]:
		  /**/
		  (r_counter==200) ? i_data[15:0]:
		  /**/
		  (r_counter==201) ? i_data[15:0]:
		  /**/
		  (r_counter==202) ? i_data[15:0]:
		  /**/
		  (r_counter==203) ? i_data[15:0]:
		  /**/
		  (r_counter==204) ? i_data[15:0]:
		  /**/
		  (r_counter==205) ? i_data[15:0]:
		  /**/
		  (r_counter==206) ? i_data[15:0]:
		  /**/
		  (r_counter==207) ? i_data[15:0]:
		  /**/
		  (r_counter==208) ? i_data[15:0]:
		  /**/
		  (r_counter==209) ? i_data[15:0]:
		  /**/
		  (r_counter==210) ? i_data[15:0]:
		  /**/
		  (r_counter==211) ? i_data[15:0]:
		  /**/
		  (r_counter==212) ? i_data[15:0]:
		  /**/
		  (r_counter==213) ? i_data[15:0]:
		  /**/
		  (r_counter==214) ? i_data[15:0]:
		  /**/
		  (r_counter==215) ? i_data[15:0]:
		  /**/
		  (r_counter==216) ? i_data[15:0]:
		  /**/
		  (r_counter==217) ? i_data[15:0]:
		  /**/
		  (r_counter==218) ? i_data[15:0]:
		  /**/
		  (r_counter==219) ? i_data[15:0]:
		  /**/
		  (r_counter==220) ? i_data[15:0]:
		  /**/
		  (r_counter==221) ? i_data[15:0]:
		  /**/
		  (r_counter==222) ? i_data[15:0]:
		  /**/
		  (r_counter==223) ? i_data[15:0]:
		  /**/
		  (r_counter==224) ? i_data[15:0]:
		  /**/
		  (r_counter==225) ? i_data[15:0]:
		  /**/
		  (r_counter==226) ? i_data[15:0]:
		  /**/
		  (r_counter==227) ? i_data[15:0]:
		  /**/
		  (r_counter==228) ? i_data[15:0]:
		  /**/
		  (r_counter==229) ? i_data[15:0]:
		  /**/
		  (r_counter==230) ? i_data[15:0]:
		  /**/
		  (r_counter==231) ? i_data[15:0]:
		  /**/
		  (r_counter==232) ? i_data[15:0]:
		  /**/
		  (r_counter==233) ? i_data[15:0]:
		  /**/
		  (r_counter==234) ? i_data[15:0]:
		  /**/
		  (r_counter==235) ? i_data[15:0]:
		  /**/
		  (r_counter==236) ? i_data[15:0]:
		  /**/
		  (r_counter==237) ? i_data[15:0]:
		  /**/
		  (r_counter==238) ? i_data[15:0]:
		  /**/
		  (r_counter==239) ? i_data[15:0]:
		  /**/
		  (r_counter==240) ? i_data[15:0]:
		  /**/
		  (r_counter==241) ? i_data[15:0]:
		  /**/
		  (r_counter==242) ? i_data[15:0]:
		  /**/
		  (r_counter==243) ? i_data[15:0]:
		  /**/
		  (r_counter==244) ? i_data[15:0]:
		  /**/
		  (r_counter==245) ? i_data[15:0]:
		  /**/
		  (r_counter==246) ? i_data[15:0]:
		  /**/
		  (r_counter==247) ? i_data[15:0]:
		  /**/
		  (r_counter==248) ? i_data[15:0]:
		  /**/
		  (r_counter==249) ? i_data[15:0]:
		  /**/
		  (r_counter==250) ? i_data[15:0]:
		  /**/
		  (r_counter==251) ? i_data[15:0]:
		  /**/
		  (r_counter==252) ? i_data[15:0]:
		  /**/
		  (r_counter==253) ? i_data[15:0]:
		  /**/
		  (r_counter==254) ? i_data[15:0]:
		  /**/
		  (r_counter==255) ? i_data[15:0]:
		  /**/
		  (r_counter==256) ? i_data[15:0]:
		  /**/
		  (r_counter==257) ? i_data[15:0]:
		  /**/
		  (r_counter==258) ? i_data[15:0]:
		  /**/
		  (r_counter==259) ? i_data[15:0]:
		  /**/
		  (r_counter==260) ? i_data[15:0]:
		  /**/
		  (r_counter==261) ? i_data[15:0]:
		  /**/
		  (r_counter==262) ? i_data[15:0]:
		  /**/
		  (r_counter==263) ? i_data[15:0]:
		  /**/
		  (r_counter==264) ? i_data[15:0]:
		  /**/
		  (r_counter==265) ? i_data[15:0]:
		  /**/
		  (r_counter==266) ? i_data[15:0]:
		  /**/
		  (r_counter==267) ? i_data[15:0]:
		  /**/
		  (r_counter==268) ? i_data[15:0]:
		  /**/
		  (r_counter==269) ? i_data[15:0]:
		  /**/
		  (r_counter==270) ? i_data[15:0]:
		  /**/
		  (r_counter==271) ? i_data[15:0]:
		  /**/
		  (r_counter==272) ? i_data[15:0]:
		  /**/
		  (r_counter==273) ? i_data[15:0]:
		  /**/
		  (r_counter==274) ? i_data[15:0]:
		  /**/
		  (r_counter==275) ? i_data[15:0]:
		  /**/
		  (r_counter==276) ? i_data[15:0]:
		  /**/
		  (r_counter==277) ? i_data[15:0]:
		  /**/
		  (r_counter==278) ? i_data[15:0]:
		  /**/
		  (r_counter==279) ? i_data[15:0]:
		  /**/
		  (r_counter==280) ? i_data[15:0]:
		  /**/
		  (r_counter==281) ? i_data[15:0]:
		  /**/
		  (r_counter==282) ? i_data[15:0]:
		  /**/
		  (r_counter==283) ? i_data[15:0]:
		  /**/
		  (r_counter==284) ? i_data[15:0]:
		  /**/
		  (r_counter==285) ? i_data[15:0]:
		  /**/
		  (r_counter==286) ? i_data[15:0]:
		  /**/
		  (r_counter==287) ? i_data[15:0]:
		  /**/
		  (r_counter==288) ? i_data[15:0]:
		  /**/
		  (r_counter==289) ? i_data[15:0]:
		  /**/
		  (r_counter==290) ? i_data[15:0]:
		  /**/
		  (r_counter==291) ? i_data[15:0]:
		  /**/
		  (r_counter==292) ? i_data[15:0]:
		  /**/
		  (r_counter==293) ? i_data[15:0]:
		  /**/
		  (r_counter==294) ? i_data[15:0]:
		  /**/
		  (r_counter==295) ? i_data[15:0]:
		  /**/
		  (r_counter==296) ? i_data[15:0]:
		  /**/
		  (r_counter==297) ? i_data[15:0]:
		  /**/
		  (r_counter==298) ? i_data[15:0]:
		  /**/
		  (r_counter==299) ? i_data[15:0]:
		  /**/
		  (r_counter==300) ? i_data[15:0]:
		  /**/
		  (r_counter==301) ? i_data[15:0]:
		  /**/
		  (r_counter==302) ? i_data[15:0]:
		  /**/
		  (r_counter==303) ? i_data[15:0]:
		  /**/
		  (r_counter==304) ? i_data[15:0]:
		  /**/
		  (r_counter==305) ? i_data[15:0]:
		  /**/
		  (r_counter==306) ? i_data[15:0]:
		  /**/
		  (r_counter==307) ? i_data[15:0]:
		  /**/
		  (r_counter==308) ? i_data[15:0]:
		  /**/
		  (r_counter==309) ? i_data[15:0]:
		  /**/
		  (r_counter==310) ? i_data[15:0]:
		  /**/
		  (r_counter==311) ? i_data[15:0]:
		  /**/
		  (r_counter==312) ? i_data[15:0]:
		  /**/
		  (r_counter==313) ? i_data[15:0]:
		  /**/
		  (r_counter==314) ? i_data[15:0]:
		  /**/
		  (r_counter==315) ? i_data[15:0]:
		  /**/
		  (r_counter==316) ? i_data[15:0]:
		  /**/
		  (r_counter==317) ? i_data[15:0]:
		  /**/
		  (r_counter==318) ? i_data[15:0]:
		  /**/
		  (r_counter==319) ? i_data[15:0]:
		  /**/
		  (r_counter==320) ? i_data[15:0]:
		  /**/
		  (r_counter==321) ? i_data[15:0]:
		  /**/
		  (r_counter==322) ? i_data[15:0]:
		  /**/
		  (r_counter==323) ? i_data[15:0]:
		  /**/
		  (r_counter==324) ? i_data[15:0]:
		  /**/
		  (r_counter==325) ? i_data[15:0]:
		  /**/
		  (r_counter==326) ? i_data[15:0]:
		  /**/
		  (r_counter==327) ? i_data[15:0]:
		  /**/
		  (r_counter==328) ? i_data[15:0]:
		  /**/
		  (r_counter==329) ? i_data[15:0]:
		  /**/
		  (r_counter==330) ? i_data[15:0]:
		  /**/
		  (r_counter==331) ? i_data[15:0]:
		  /**/
		  (r_counter==332) ? i_data[15:0]:
		  /**/
		  (r_counter==333) ? i_data[15:0]:
		  /**/
		  (r_counter==334) ? i_data[15:0]:
		  /**/
		  (r_counter==335) ? i_data[15:0]:
		  /**/
		  (r_counter==336) ? i_data[15:0]:
		  /**/
		  (r_counter==337) ? i_data[15:0]:
		  /**/
		  (r_counter==338) ? i_data[15:0]:
		  /**/
		  (r_counter==339) ? i_data[15:0]:
		  /**/
		  (r_counter==340) ? i_data[15:0]:
		  /**/
		  (r_counter==341) ? i_data[15:0]:
		  /**/
		  (r_counter==342) ? i_data[15:0]:
		  /**/
		  (r_counter==343) ? i_data[15:0]:
		  /**/
		  (r_counter==344) ? i_data[15:0]:
		  /**/
		  (r_counter==345) ? i_data[15:0]:
		  /**/
		  (r_counter==346) ? i_data[15:0]:
		  /**/
		  (r_counter==347) ? i_data[15:0]:
		  /**/
		  (r_counter==348) ? i_data[15:0]:
		  /**/
		  (r_counter==349) ? i_data[15:0]:
		  /**/
		  (r_counter==350) ? i_data[15:0]:
		  /**/
		  (r_counter==351) ? i_data[15:0]:
		  /**/
		  (r_counter==352) ? i_data[15:0]:
		  /**/
		  (r_counter==353) ? i_data[15:0]:
		  /**/
		  (r_counter==354) ? i_data[15:0]:
		  /**/
		  (r_counter==355) ? i_data[15:0]:
		  /**/
		  (r_counter==356) ? i_data[15:0]:
		  /**/
		  (r_counter==357) ? i_data[15:0]:
		  /**/
		  (r_counter==358) ? i_data[15:0]:
		  /**/
		  (r_counter==359) ? i_data[15:0]:
		  /**/
		  (r_counter==360) ? i_data[15:0]:
		  /**/
		  (r_counter==361) ? i_data[15:0]:
		  /**/
		  (r_counter==362) ? i_data[15:0]:
		  /**/
		  (r_counter==363) ? i_data[15:0]:
		  /**/
		  (r_counter==364) ? i_data[15:0]:
		  /**/
		  (r_counter==365) ? i_data[15:0]:
		  /**/
		  (r_counter==366) ? i_data[15:0]:
		  /**/
		  (r_counter==367) ? i_data[15:0]:
		  /**/
		  (r_counter==368) ? i_data[15:0]:
		  /**/
		  (r_counter==369) ? i_data[15:0]:
		  /**/
		  (r_counter==370) ? i_data[15:0]:
		  /**/
		  (r_counter==371) ? i_data[15:0]:
		  /**/
		  (r_counter==372) ? i_data[15:0]:
		  /**/
		  (r_counter==373) ? i_data[15:0]:
		  /**/
		  (r_counter==374) ? i_data[15:0]:
		  /**/
		  (r_counter==375) ? i_data[15:0]:
		  /**/
		  (r_counter==376) ? i_data[15:0]:
		  /**/
		  (r_counter==377) ? i_data[15:0]:
		  /**/
		  (r_counter==378) ? i_data[15:0]:
		  /**/
		  (r_counter==379) ? i_data[15:0]:
		  /**/
		  (r_counter==380) ? i_data[15:0]:
		  /**/
		  (r_counter==381) ? i_data[15:0]:
		  /**/
		  (r_counter==382) ? i_data[15:0]:
		  /**/
		  (r_counter==383) ? i_data[15:0]:
		  /**/
		  (r_counter==384) ? i_data[15:0]:
		  /**/
		  (r_counter==385) ? i_data[15:0]:
		  /**/
		  (r_counter==386) ? i_data[15:0]:
		  /**/
		  (r_counter==387) ? i_data[15:0]:
		  /**/
		  (r_counter==388) ? i_data[15:0]:
		  /**/
		  (r_counter==389) ? i_data[15:0]:
		  /**/
		  (r_counter==390) ? i_data[15:0]:
		  /**/
		  (r_counter==391) ? i_data[15:0]:
		  /**/
		  (r_counter==392) ? i_data[15:0]:
		  /**/
		  (r_counter==393) ? i_data[15:0]:
		  /**/
		  (r_counter==394) ? i_data[15:0]:
		  /**/
		  (r_counter==395) ? i_data[15:0]:
		  /**/
		  (r_counter==396) ? i_data[15:0]:
		  /**/
		  (r_counter==397) ? i_data[15:0]:
		  /**/
		  (r_counter==398) ? i_data[15:0]:
		  /**/
		  (r_counter==399) ? i_data[15:0]:
		  /**/
		  0;
   //alpha
   assign i_wen_alpha=(r_state==zStateRow) & (
					      /**/
					      (r_counter == (4)) |
					      /**/
					      (r_counter == (7)) |
					      /**/
					      (r_counter == (10)) |
					      /**/
					      (r_counter == (13)) |
					      /**/
					      (r_counter == (16)) |
					      /**/
					      (r_counter == (19)) |
					      /**/
					      (r_counter == (22)) |
					      /**/
					      (r_counter == (25)) |
					      /**/
					      (r_counter == (28)) |
					      /**/
					      (r_counter == (31)) |
					      /**/
					      (r_counter == (34)) |
					      /**/
					      (r_counter == (37)) |
					      /**/
					      (r_counter == (40)) |
					      /**/
					      (r_counter == (43)) |
					      /**/
					      (r_counter == (46)) |
					      /**/
					      (r_counter == (49)) |
					      /**/
					      (r_counter == (52)) |
					      /**/
					      (r_counter == (55)) |
					      /**/
					      (r_counter == (58)) |
					      /**/
					      (r_counter == (61)) |
					      /**/
					      (r_counter == (64)) |
					      /**/
					      (r_counter == (67)) |
					      /**/
					      (r_counter == (70)) |
					      /**/
					      (r_counter == (73)) |
					      /**/
					      (r_counter == (76)) |
					      /**/
					      (r_counter == (79)) |
					      /**/
					      (r_counter == (82)) |
					      /**/
					      (r_counter == (85)) |
					      /**/
					      (r_counter == (88)) |
					      /**/
					      (r_counter == (91)) |
					      /**/
					      (r_counter == (94)) |
					      /**/
					      (r_counter == (97)) |
					      /**/
					      (r_counter == (100)) |
					      /**/
					      (r_counter == (103)) |
					      /**/
					      (r_counter == (106)) |
					      /**/
					      (r_counter == (109)) |
					      /**/
					      (r_counter == (112)) |
					      /**/
					      (r_counter == (115)) |
					      /**/
					      (r_counter == (118)) |
					      /**/
					      (r_counter == (121)) |
					      /**/
					      (r_counter == (124)) |
					      /**/
					      (r_counter == (127)) |
					      /**/
					      (r_counter == (130)) |
					      /**/
					      (r_counter == (133)) |
					      /**/
					      (r_counter == (136)) |
					      /**/
					      (r_counter == (139)) |
					      /**/
					      (r_counter == (142)) |
					      /**/
					      (r_counter == (145)) |
					      /**/
					      (r_counter == (148)) |
					      /**/
					      (r_counter == (151)) |
					      /**/
					      (r_counter == (154)) |
					      /**/
					      (r_counter == (157)) |
					      /**/
					      (r_counter == (160)) |
					      /**/
					      (r_counter == (163)) |
					      /**/
					      (r_counter == (166)) |
					      /**/
					      (r_counter == (169)) |
					      /**/
					      (r_counter == (172)) |
					      /**/
					      (r_counter == (175)) |
					      /**/
					      (r_counter == (178)) |
					      /**/
					      (r_counter == (181)) |
					      /**/
					      (r_counter == (184)) |
					      /**/
					      (r_counter == (187)) |
					      /**/
					      (r_counter == (190)) |
					      /**/
					      (r_counter == (193)) |
					      /**/
					      (r_counter == (196)) |
					      /**/
					      (r_counter == (199)) |
					      /**/
					      (r_counter == (202)) |
					      /**/
					      (r_counter == (205)) |
					      /**/
					      (r_counter == (208)) |
					      /**/
					      (r_counter == (211)) |
					      /**/
					      (r_counter == (214)) |
					      /**/
					      (r_counter == (217)) |
					      /**/
					      (r_counter == (220)) |
					      /**/
					      (r_counter == (223)) |
					      /**/
					      (r_counter == (226)) |
					      /**/
					      (r_counter == (229)) |
					      /**/
					      (r_counter == (232)) |
					      /**/
					      (r_counter == (235)) |
					      /**/
					      (r_counter == (238)) |
					      /**/
					      (r_counter == (241)) |
					      /**/
					      (r_counter == (244)) |
					      /**/
					      (r_counter == (247)) |
					      /**/
					      (r_counter == (250)) |
					      /**/
					      (r_counter == (253)) |
					      /**/
					      (r_counter == (256)) |
					      /**/
					      (r_counter == (259)) |
					      /**/
					      (r_counter == (262)) |
					      /**/
					      (r_counter == (265)) |
					      /**/
					      (r_counter == (268)) |
					      /**/
					      (r_counter == (271)) |
					      /**/
					      (r_counter == (274)) |
					      /**/
					      (r_counter == (277)) |
					      /**/
					      (r_counter == (280)) |
					      /**/
					      (r_counter == (283)) |
					      /**/
					      (r_counter == (286)) |
					      /**/
					      (r_counter == (289)) |
					      /**/
					      (r_counter == (292)) |
					      /**/
					      (r_counter == (295)) |
					      /**/
					      (r_counter == (298)) |
					      /**/
					      (r_counter == (301)) |
					      /**/
					      (r_counter == (304)) |
					      /**/
					      (r_counter == (307)) |
					      /**/
					      (r_counter == (310)) |
					      /**/
					      (r_counter == (313)) |
					      /**/
					      (r_counter == (316)) |
					      /**/
					      (r_counter == (319)) |
					      /**/
					      (r_counter == (322)) |
					      /**/
					      (r_counter == (325)) |
					      /**/
					      (r_counter == (328)) |
					      /**/
					      (r_counter == (331)) |
					      /**/
					      (r_counter == (334)) |
					      /**/
					      (r_counter == (337)) |
					      /**/
					      (r_counter == (340)) |
					      /**/
					      (r_counter == (343)) |
					      /**/
					      (r_counter == (346)) |
					      /**/
					      (r_counter == (349)) |
					      /**/
					      (r_counter == (352)) |
					      /**/
					      (r_counter == (355)) |
					      /**/
					      (r_counter == (358)) |
					      /**/
					      (r_counter == (361)) |
					      /**/
					      (r_counter == (364)) |
					      /**/
					      (r_counter == (367)) |
					      /**/
					      (r_counter == (370)) |
					      /**/
					      (r_counter == (373)) |
					      /**/
					      (r_counter == (376)) |
					      /**/
					      (r_counter == (379)) |
					      /**/
					      (r_counter == (382)) |
					      /**/
					      (r_counter == (385)) |
					      /**/
					      (r_counter == (388)) |
					      /**/
					      (r_counter == (391)) |
					      /**/
					      (r_counter == (394)) |
					      /**/
					      (r_counter == (397)) |
					      /**/
					      (r_counter == (400)) |
					      /**/
					      (r_counter == (403)) |
					      /**/
					      (r_counter == (406)) |
					      /**/
					      (r_counter == (409)) |
					      /**/
					      (r_counter == (412)) |
					      /**/
					      (r_counter == (415)) |
					      /**/
					      (r_counter == (418)) |
					      /**/
					      (r_counter == (421)) |
					      /**/
					      (r_counter == (424)) |
					      /**/
					      (r_counter == (427)) |
					      /**/
					      (r_counter == (430)) |
					      /**/
					      (r_counter == (433)) |
					      /**/
					      (r_counter == (436)) |
					      /**/
					      (r_counter == (439)) |
					      /**/
					      (r_counter == (442)) |
					      /**/
					      (r_counter == (445)) |
					      /**/
					      (r_counter == (448)) |
					      /**/
					      (r_counter == (451)) |
					      /**/
					      (r_counter == (454)) |
					      /**/
					      (r_counter == (457)) |
					      /**/
					      (r_counter == (460)) |
					      /**/
					      (r_counter == (463)) |
					      /**/
					      (r_counter == (466)) |
					      /**/
					      (r_counter == (469)) |
					      /**/
					      (r_counter == (472)) |
					      /**/
					      (r_counter == (475)) |
					      /**/
					      (r_counter == (478)) |
					      /**/
					      (r_counter == (481)) |
					      /**/
					      (r_counter == (484)) |
					      /**/
					      (r_counter == (487)) |
					      /**/
					      (r_counter == (490)) |
					      /**/
					      (r_counter == (493)) |
					      /**/
					      (r_counter == (496)) |
					      /**/
					      (r_counter == (499)) |
					      /**/
					      (r_counter == (502)) |
					      /**/
					      (r_counter == (505)) |
					      /**/
					      (r_counter == (508)) |
					      /**/
					      (r_counter == (511)) |
					      /**/
					      (r_counter == (514)) |
					      /**/
					      (r_counter == (517)) |
					      /**/
					      (r_counter == (520)) |
					      /**/
					      (r_counter == (523)) |
					      /**/
					      (r_counter == (526)) |
					      /**/
					      (r_counter == (529)) |
					      /**/
					      (r_counter == (532)) |
					      /**/
					      (r_counter == (535)) |
					      /**/
					      (r_counter == (538)) |
					      /**/
					      (r_counter == (541)) |
					      /**/
					      (r_counter == (544)) |
					      /**/
					      (r_counter == (547)) |
					      /**/
					      (r_counter == (550)) |
					      /**/
					      (r_counter == (553)) |
					      /**/
					      (r_counter == (556)) |
					      /**/
					      (r_counter == (559)) |
					      /**/
					      (r_counter == (562)) |
					      /**/
					      (r_counter == (565)) |
					      /**/
					      (r_counter == (568)) |
					      /**/
					      (r_counter == (571)) |
					      /**/
					      (r_counter == (574)) |
					      /**/
					      (r_counter == (577)) |
					      /**/
					      (r_counter == (580)) |
					      /**/
					      (r_counter == (583)) |
					      /**/
					      (r_counter == (586)) |
					      /**/
					      (r_counter == (589)) |
					      /**/
					      (r_counter == (592)) |
					      /**/
					      (r_counter == (595)) |
					      /**/
					      (r_counter == (598)) |
					      /**/
					      (r_counter == (601)) |
					      /**/
					      (r_counter == (604)) |
					      /**/
					      (r_counter == (607)) |
					      /**/
					      (r_counter == (610)) |
					      /**/
					      (r_counter == (613)) |
					      /**/
					      (r_counter == (616)) |
					      /**/
					      (r_counter == (619)) |
					      /**/
					      (r_counter == (622)) |
					      /**/
					      (r_counter == (625)) |
					      /**/
					      (r_counter == (628)) |
					      /**/
					      (r_counter == (631)) |
					      /**/
					      (r_counter == (634)) |
					      /**/
					      (r_counter == (637)) |
					      /**/
					      (r_counter == (640)) |
					      /**/
					      (r_counter == (643)) |
					      /**/
					      (r_counter == (646)) |
					      /**/
					      (r_counter == (649)) |
					      /**/
					      (r_counter == (652)) |
					      /**/
					      (r_counter == (655)) |
					      /**/
					      (r_counter == (658)) |
					      /**/
					      (r_counter == (661)) |
					      /**/
					      (r_counter == (664)) |
					      /**/
					      (r_counter == (667)) |
					      /**/
					      (r_counter == (670)) |
					      /**/
					      (r_counter == (673)) |
					      /**/
					      (r_counter == (676)) |
					      /**/
					      (r_counter == (679)) |
					      /**/
					      (r_counter == (682)) |
					      /**/
					      (r_counter == (685)) |
					      /**/
					      (r_counter == (688)) |
					      /**/
					      (r_counter == (691)) |
					      /**/
					      (r_counter == (694)) |
					      /**/
					      (r_counter == (697)) |
					      /**/
					      (r_counter == (700)) |
					      /**/
					      (r_counter == (703)) |
					      /**/
					      (r_counter == (706)) |
					      /**/
					      (r_counter == (709)) |
					      /**/
					      (r_counter == (712)) |
					      /**/
					      (r_counter == (715)) |
					      /**/
					      (r_counter == (718)) |
					      /**/
					      (r_counter == (721)) |
					      /**/
					      (r_counter == (724)) |
					      /**/
					      (r_counter == (727)) |
					      /**/
					      (r_counter == (730)) |
					      /**/
					      (r_counter == (733)) |
					      /**/
					      (r_counter == (736)) |
					      /**/
					      (r_counter == (739)) |
					      /**/
					      (r_counter == (742)) |
					      /**/
					      (r_counter == (745)) |
					      /**/
					      (r_counter == (748)) |
					      /**/
					      (r_counter == (751)) |
					      /**/
					      (r_counter == (754)) |
					      /**/
					      (r_counter == (757)) |
					      /**/
					      (r_counter == (760)) |
					      /**/
					      (r_counter == (763)) |
					      /**/
					      (r_counter == (766)) |
					      /**/
					      (r_counter == (769)) |
					      /**/
					      (r_counter == (772)) |
					      /**/
					      (r_counter == (775)) |
					      /**/
					      (r_counter == (778)) |
					      /**/
					      (r_counter == (781)) |
					      /**/
					      (r_counter == (784)) |
					      /**/
					      (r_counter == (787)) |
					      /**/
					      (r_counter == (790)) |
					      /**/
					      (r_counter == (793)) |
					      /**/
					      (r_counter == (796)) |
					      /**/
					      (r_counter == (799)) |
					      /**/
					      (r_counter == (802)) |
					      /**/
					      (r_counter == (805)) |
					      /**/
					      (r_counter == (808)) |
					      /**/
					      (r_counter == (811)) |
					      /**/
					      (r_counter == (814)) |
					      /**/
					      (r_counter == (817)) |
					      /**/
					      (r_counter == (820)) |
					      /**/
					      (r_counter == (823)) |
					      /**/
					      (r_counter == (826)) |
					      /**/
					      (r_counter == (829)) |
					      /**/
					      (r_counter == (832)) |
					      /**/
					      (r_counter == (835)) |
					      /**/
					      (r_counter == (838)) |
					      /**/
					      (r_counter == (841)) |
					      /**/
					      (r_counter == (844)) |
					      /**/
					      (r_counter == (847)) |
					      /**/
					      (r_counter == (850)) |
					      /**/
					      (r_counter == (853)) |
					      /**/
					      (r_counter == (856)) |
					      /**/
					      (r_counter == (859)) |
					      /**/
					      (r_counter == (862)) |
					      /**/
					      (r_counter == (865)) |
					      /**/
					      (r_counter == (868)) |
					      /**/
					      (r_counter == (871)) |
					      /**/
					      (r_counter == (874)) |
					      /**/
					      (r_counter == (877)) |
					      /**/
					      (r_counter == (880)) |
					      /**/
					      (r_counter == (883)) |
					      /**/
					      (r_counter == (886)) |
					      /**/
					      (r_counter == (889)) |
					      /**/
					      (r_counter == (892)) |
					      /**/
					      (r_counter == (895)) |
					      /**/
					      (r_counter == (898)) |
					      /**/
					      (r_counter == (901)) |
					      /**/
					      (r_counter == (904)) |
					      /**/
					      (r_counter == (907)) |
					      /**/
					      (r_counter == (910)) |
					      /**/
					      (r_counter == (913)) |
					      /**/
					      (r_counter == (916)) |
					      /**/
					      (r_counter == (919)) |
					      /**/
					      (r_counter == (922)) |
					      /**/
					      (r_counter == (925)) |
					      /**/
					      (r_counter == (928)) |
					      /**/
					      (r_counter == (931)) |
					      /**/
					      (r_counter == (934)) |
					      /**/
					      (r_counter == (937)) |
					      /**/
					      (r_counter == (940)) |
					      /**/
					      (r_counter == (943)) |
					      /**/
					      (r_counter == (946)) |
					      /**/
					      (r_counter == (949)) |
					      /**/
					      (r_counter == (952)) |
					      /**/
					      (r_counter == (955)) |
					      /**/
					      (r_counter == (958)) |
					      /**/
					      (r_counter == (961)) |
					      /**/
					      (r_counter == (964)) |
					      /**/
					      (r_counter == (967)) |
					      /**/
					      (r_counter == (970)) |
					      /**/
					      (r_counter == (973)) |
					      /**/
					      (r_counter == (976)) |
					      /**/
					      (r_counter == (979)) |
					      /**/
					      (r_counter == (982)) |
					      /**/
					      (r_counter == (985)) |
					      /**/
					      (r_counter == (988)) |
					      /**/
					      (r_counter == (991)) |
					      /**/
					      (r_counter == (994)) |
					      /**/
					      (r_counter == (997)) |
					      /**/
					      (r_counter == (1000)) |
					      /**/
					      (r_counter == (1003)) |
					      /**/
					      (r_counter == (1006)) |
					      /**/
					      (r_counter == (1009)) |
					      /**/
					      (r_counter == (1012)) |
					      /**/
					      (r_counter == (1015)) |
					      /**/
					      (r_counter == (1018)) |
					      /**/
					      (r_counter == (1021)) |
					      /**/
					      (r_counter == (1024)) |
					      /**/
					      (r_counter == (1027)) |
					      /**/
					      (r_counter == (1030)) |
					      /**/
					      (r_counter == (1033)) |
					      /**/
					      (r_counter == (1036)) |
					      /**/
					      (r_counter == (1039)) |
					      /**/
					      (r_counter == (1042)) |
					      /**/
					      (r_counter == (1045)) |
					      /**/
					      (r_counter == (1048)) |
					      /**/
					      (r_counter == (1051)) |
					      /**/
					      (r_counter == (1054)) |
					      /**/
					      (r_counter == (1057)) |
					      /**/
					      (r_counter == (1060)) |
					      /**/
					      (r_counter == (1063)) |
					      /**/
					      (r_counter == (1066)) |
					      /**/
					      (r_counter == (1069)) |
					      /**/
					      (r_counter == (1072)) |
					      /**/
					      (r_counter == (1075)) |
					      /**/
					      (r_counter == (1078)) |
					      /**/
					      (r_counter == (1081)) |
					      /**/
					      (r_counter == (1084)) |
					      /**/
					      (r_counter == (1087)) |
					      /**/
					      (r_counter == (1090)) |
					      /**/
					      (r_counter == (1093)) |
					      /**/
					      (r_counter == (1096)) |
					      /**/
					      (r_counter == (1099)) |
					      /**/
					      (r_counter == (1102)) |
					      /**/
					      (r_counter == (1105)) |
					      /**/
					      (r_counter == (1108)) |
					      /**/
					      (r_counter == (1111)) |
					      /**/
					      (r_counter == (1114)) |
					      /**/
					      (r_counter == (1117)) |
					      /**/
					      (r_counter == (1120)) |
					      /**/
					      (r_counter == (1123)) |
					      /**/
					      (r_counter == (1126)) |
					      /**/
					      (r_counter == (1129)) |
					      /**/
					      (r_counter == (1132)) |
					      /**/
					      (r_counter == (1135)) |
					      /**/
					      (r_counter == (1138)) |
					      /**/
					      (r_counter == (1141)) |
					      /**/
					      (r_counter == (1144)) |
					      /**/
					      (r_counter == (1147)) |
					      /**/
					      (r_counter == (1150)) |
					      /**/
					      (r_counter == (1153)) |
					      /**/
					      (r_counter == (1156)) |
					      /**/
					      (r_counter == (1159)) |
					      /**/
					      (r_counter == (1162)) |
					      /**/
					      (r_counter == (1165)) |
					      /**/
					      (r_counter == (1168)) |
					      /**/
					      (r_counter == (1171)) |
					      /**/
					      (r_counter == (1174)) |
					      /**/
					      (r_counter == (1177)) |
					      /**/
					      (r_counter == (1180)) |
					      /**/
					      (r_counter == (1183)) |
					      /**/
					      (r_counter == (1186)) |
					      /**/
					      (r_counter == (1189)) |
					      /**/
					      (r_counter == (1192)) |
					      /**/
					      (r_counter == (1195)) |
					      /**/
					      (r_counter == (1198)) |
					      /**/
					      (r_counter == (1201)) |
					      /**/
					      (r_counter == (1204)) |
					      /**/
					      (r_counter == (1207)) |
					      /**/
					      (r_counter == (1210)) |
					      /**/
					      (r_counter == (1213)) |
					      /**/
					      (r_counter == (1216)) |
					      /**/
					      (r_counter == (1219)) |
					      /**/
					      (r_counter == (1222)) |
					      /**/
					      (r_counter == (1225)) |
					      /**/
					      (r_counter == (1228)) |
					      /**/
					      (r_counter == (1231)) |
					      /**/
					      (r_counter == (1234)) |
					      /**/
					      (r_counter == (1237)) |
					      /**/
					      (r_counter == (1240)) |
					      /**/
					      (r_counter == (1243)) |
					      /**/
					      (r_counter == (1246)) |
					      /**/
					      (r_counter == (1249)) |
					      /**/
					      (r_counter == (1252)) |
					      /**/
					      (r_counter == (1255)) |
					      /**/
					      (r_counter == (1258)) |
					      /**/
					      (r_counter == (1261)) |
					      /**/
					      (r_counter == (1264)) |
					      /**/
					      (r_counter == (1267)) |
					      /**/
					      (r_counter == (1270)) |
					      /**/
					      (r_counter == (1273)) |
					      /**/
					      (r_counter == (1276)) |
					      /**/
					      (r_counter == (1279)) |
					      /**/
					      (r_counter == (1282)) |
					      /**/
					      (r_counter == (1285)) |
					      /**/
					      (r_counter == (1288)) |
					      /**/
					      (r_counter == (1291)) |
					      /**/
					      (r_counter == (1294)) |
					      /**/
					      (r_counter == (1297)) |
					      /**/
					      (r_counter == (1300)) |
					      /**/
					      (r_counter == (1303)) |
					      /**/
					      (r_counter == (1306)) |
					      /**/
					      (r_counter == (1309)) |
					      /**/
					      (r_counter == (1312)) |
					      /**/
					      (r_counter == (1315)) |
					      /**/
					      (r_counter == (1318)) |
					      /**/
					      (r_counter == (1321)) |
					      /**/
					      (r_counter == (1324)) |
					      /**/
					      (r_counter == (1327)) |
					      /**/
					      (r_counter == (1330)) |
					      /**/
					      (r_counter == (1333)) |
					      /**/
					      (r_counter == (1336)) |
					      /**/
					      (r_counter == (1339)) |
					      /**/
					      (r_counter == (1342)) |
					      /**/
					      (r_counter == (1345)) |
					      /**/
					      (r_counter == (1348)) |
					      /**/
					      (r_counter == (1351)) |
					      /**/
					      (r_counter == (1354)) |
					      /**/
					      (r_counter == (1357)) |
					      /**/
					      (r_counter == (1360)) |
					      /**/
					      (r_counter == (1363)) |
					      /**/
					      (r_counter == (1366)) |
					      /**/
					      (r_counter == (1369)) |
					      /**/
					      (r_counter == (1372)) |
					      /**/
					      (r_counter == (1375)) |
					      /**/
					      (r_counter == (1378)) |
					      /**/
					      (r_counter == (1381)) |
					      /**/
					      (r_counter == (1384)) |
					      /**/
					      (r_counter == (1387)) |
					      /**/
					      (r_counter == (1390)) |
					      /**/
					      (r_counter == (1393)) |
					      /**/
					      (r_counter == (1396)) |
					      /**/
					      (r_counter == (1399)) |
					      /**/
					      (r_counter == (1402)) |
					      /**/
					      (r_counter == (1405)) |
					      /**/
					      (r_counter == (1408)) |
					      /**/
					      (r_counter == (1411)) |
					      /**/
					      (r_counter == (1414)) |
					      /**/
					      (r_counter == (1417)) |
					      /**/
					      (r_counter == (1420)) |
					      /**/
					      (r_counter == (1423)) |
					      /**/
					      (r_counter == (1426)) |
					      /**/
					      (r_counter == (1429)) |
					      /**/
					      (r_counter == (1432)) |
					      /**/
					      (r_counter == (1435)) |
					      /**/
					      (r_counter == (1438)) |
					      /**/
					      (r_counter == (1441)) |
					      /**/
					      (r_counter == (1444)) |
					      /**/
					      (r_counter == (1447)) |
					      /**/
					      (r_counter == (1450)) |
					      /**/
					      (r_counter == (1453)) |
					      /**/
					      (r_counter == (1456)) |
					      /**/
					      (r_counter == (1459)) |
					      /**/
					      (r_counter == (1462)) |
					      /**/
					      (r_counter == (1465)) |
					      /**/
					      (r_counter == (1468)) |
					      /**/
					      (r_counter == (1471)) |
					      /**/
					      (r_counter == (1474)) |
					      /**/
					      (r_counter == (1477)) |
					      /**/
					      (r_counter == (1480)) |
					      /**/
					      (r_counter == (1483)) |
					      /**/
					      (r_counter == (1486)) |
					      /**/
					      (r_counter == (1489)) |
					      /**/
					      (r_counter == (1492)) |
					      /**/
					      (r_counter == (1495)) |
					      /**/
					      (r_counter == (1498)) |
					      /**/
					      (r_counter == (1501)) |
					      /**/
					      (r_counter == (1504)) |
					      /**/
					      (r_counter == (1507)) |
					      /**/
					      (r_counter == (1510)) |
					      /**/
					      (r_counter == (1513)) |
					      /**/
					      (r_counter == (1516)) |
					      /**/
					      (r_counter == (1519)) |
					      /**/
					      (r_counter == (1522)) |
					      /**/
					      (r_counter == (1525)) |
					      /**/
					      (r_counter == (1528)) |
					      /**/
					      (r_counter == (1531)) |
					      /**/
					      (r_counter == (1534)) |
					      /**/
					      (r_counter == (1537)) |
					      /**/
					      (r_counter == (1540)) |
					      /**/
					      (r_counter == (1543)) |
					      /**/
					      (r_counter == (1546)) |
					      /**/
					      (r_counter == (1549)) |
					      /**/
					      (r_counter == (1552)) |
					      /**/
					      (r_counter == (1555)) |
					      /**/
					      (r_counter == (1558)) |
					      /**/
					      (r_counter == (1561)) |
					      /**/
					      (r_counter == (1564)) |
					      /**/
					      (r_counter == (1567)) |
					      /**/
					      (r_counter == (1570)) |
					      /**/
					      (r_counter == (1573)) |
					      /**/
					      (r_counter == (1576)) |
					      /**/
					      (r_counter == (1579)) |
					      /**/
					      (r_counter == (1582)) |
					      /**/
					      (r_counter == (1585)) |
					      /**/
					      (r_counter == (1588)) |
					      /**/
					      (r_counter == (1591)) |
					      /**/
					      (r_counter == (1594)) |
					      /**/
					      (r_counter == (1597)) |
					      /**/
					      (r_counter == (1600)) |
					      /**/
					      (r_counter == (1603)) |
					      /**/
					      (r_counter == (1606)) |
					      /**/
					      (r_counter == (1609)) |
					      /**/
					      (r_counter == (1612)) |
					      /**/
					      (r_counter == (1615)) |
					      /**/
					      (r_counter == (1618)) |
					      /**/
					      (r_counter == (1621)) |
					      /**/
					      (r_counter == (1624)) |
					      /**/
					      (r_counter == (1627)) |
					      /**/
					      (r_counter == (1630)) |
					      /**/
					      (r_counter == (1633)) |
					      /**/
					      (r_counter == (1636)) |
					      /**/
					      (r_counter == (1639)) |
					      /**/
					      (r_counter == (1642)) |
					      /**/
					      (r_counter == (1645)) |
					      /**/
					      (r_counter == (1648)) |
					      /**/
					      (r_counter == (1651)) |
					      /**/
					      (r_counter == (1654)) |
					      /**/
					      (r_counter == (1657)) |
					      /**/
					      (r_counter == (1660)) |
					      /**/
					      (r_counter == (1663)) |
					      /**/
					      (r_counter == (1666)) |
					      /**/
					      (r_counter == (1669)) |
					      /**/
					      (r_counter == (1672)) |
					      /**/
					      (r_counter == (1675)) |
					      /**/
					      (r_counter == (1678)) |
					      /**/
					      (r_counter == (1681)) |
					      /**/
					      (r_counter == (1684)) |
					      /**/
					      (r_counter == (1687)) |
					      /**/
					      (r_counter == (1690)) |
					      /**/
					      (r_counter == (1693)) |
					      /**/
					      (r_counter == (1696)) |
					      /**/
					      (r_counter == (1699)) |
					      /**/
					      (r_counter == (1702)) |
					      /**/
					      (r_counter == (1705)) |
					      /**/
					      (r_counter == (1708)) |
					      /**/
					      (r_counter == (1711)) |
					      /**/
					      (r_counter == (1714)) |
					      /**/
					      (r_counter == (1717)) |
					      /**/
					      (r_counter == (1720)) |
					      /**/
					      (r_counter == (1723)) |
					      /**/
					      (r_counter == (1726)) |
					      /**/
					      (r_counter == (1729)) |
					      /**/
					      (r_counter == (1732)) |
					      /**/
					      (r_counter == (1735)) |
					      /**/
					      (r_counter == (1738)) |
					      /**/
					      (r_counter == (1741)) |
					      /**/
					      (r_counter == (1744)) |
					      /**/
					      (r_counter == (1747)) |
					      /**/
					      (r_counter == (1750)) |
					      /**/
					      (r_counter == (1753)) |
					      /**/
					      (r_counter == (1756)) |
					      /**/
					      (r_counter == (1759)) |
					      /**/
					      (r_counter == (1762)) |
					      /**/
					      (r_counter == (1765)) |
					      /**/
					      (r_counter == (1768)) |
					      /**/
					      (r_counter == (1771)) |
					      /**/
					      (r_counter == (1774)) |
					      /**/
					      (r_counter == (1777)) |
					      /**/
					      (r_counter == (1780)) |
					      /**/
					      (r_counter == (1783)) |
					      /**/
					      (r_counter == (1786)) |
					      /**/
					      (r_counter == (1789)) |
					      /**/
					      (r_counter == (1792)) |
					      /**/
					      (r_counter == (1795)) |
					      /**/
					      (r_counter == (1798)) |
					      /**/
					      (r_counter == (1801)) |
					      /**/
					      (r_counter == (1804)) |
					      /**/
					      (r_counter == (1807)) |
					      /**/
					      (r_counter == (1810)) |
					      /**/
					      (r_counter == (1813)) |
					      /**/
					      (r_counter == (1816)) |
					      /**/
					      (r_counter == (1819)) |
					      /**/
					      (r_counter == (1822)) |
					      /**/
					      (r_counter == (1825)) |
					      /**/
					      (r_counter == (1828)) |
					      /**/
					      (r_counter == (1831)) |
					      /**/
					      (r_counter == (1834)) |
					      /**/
					      (r_counter == (1837)) |
					      /**/
					      (r_counter == (1840)) |
					      /**/
					      (r_counter == (1843)) |
					      /**/
					      (r_counter == (1846)) |
					      /**/
					      (r_counter == (1849)) |
					      /**/
					      (r_counter == (1852)) |
					      /**/
					      (r_counter == (1855)) |
					      /**/
					      (r_counter == (1858)) |
					      /**/
					      (r_counter == (1861)) |
					      /**/
					      (r_counter == (1864)) |
					      /**/
					      (r_counter == (1867)) |
					      /**/
					      (r_counter == (1870)) |
					      /**/
					      (r_counter == (1873)) |
					      /**/
					      (r_counter == (1876)) |
					      /**/
					      (r_counter == (1879)) |
					      /**/
					      (r_counter == (1882)) |
					      /**/
					      (r_counter == (1885)) |
					      /**/
					      (r_counter == (1888)) |
					      /**/
					      (r_counter == (1891)) |
					      /**/
					      (r_counter == (1894)) |
					      /**/
					      (r_counter == (1897)) |
					      /**/
					      (r_counter == (1900)) |
					      /**/
					      (r_counter == (1903)) |
					      /**/
					      (r_counter == (1906)) |
					      /**/
					      (r_counter == (1909)) |
					      /**/
					      (r_counter == (1912)) |
					      /**/
					      (r_counter == (1915)) |
					      /**/
					      (r_counter == (1918)) |
					      /**/
					      (r_counter == (1921)) |
					      /**/
					      (r_counter == (1924)) |
					      /**/
					      (r_counter == (1927)) |
					      /**/
					      (r_counter == (1930)) |
					      /**/
					      (r_counter == (1933)) |
					      /**/
					      (r_counter == (1936)) |
					      /**/
					      (r_counter == (1939)) |
					      /**/
					      (r_counter == (1942)) |
					      /**/
					      (r_counter == (1945)) |
					      /**/
					      (r_counter == (1948)) |
					      /**/
					      (r_counter == (1951)) |
					      /**/
					      (r_counter == (1954)) |
					      /**/
					      (r_counter == (1957)) |
					      /**/
					      (r_counter == (1960)) |
					      /**/
					      (r_counter == (1963)) |
					      /**/
					      (r_counter == (1966)) |
					      /**/
					      (r_counter == (1969)) |
					      /**/
					      (r_counter == (1972)) |
					      /**/
					      (r_counter == (1975)) |
					      /**/
					      (r_counter == (1978)) |
					      /**/
					      (r_counter == (1981)) |
					      /**/
					      (r_counter == (1984)) |
					      /**/
					      (r_counter == (1987)) |
					      /**/
					      (r_counter == (1990)) |
					      /**/
					      (r_counter == (1993)) |
					      /**/
					      (r_counter == (1996)) |
					      /**/
					      (r_counter == (1999)) |
					      /**/
					      (r_counter == (2002)) |
					      /**/
					      (r_counter == (2005)) |
					      /**/
					      (r_counter == (2008)) |
					      /**/
					      (r_counter == (2011)) |
					      /**/
					      (r_counter == (2014)) |
					      /**/
					      (r_counter == (2017)) |
					      /**/
					      (r_counter == (2020)) |
					      /**/
					      (r_counter == (2023)) |
					      /**/
					      (r_counter == (2026)) |
					      /**/
					      (r_counter == (2029)) |
					      /**/
					      (r_counter == (2032)) |
					      /**/
					      (r_counter == (2035)) |
					      /**/
					      (r_counter == (2038)) |
					      /**/
					      (r_counter == (2041)) |
					      /**/
					      (r_counter == (2044)) |
					      /**/
					      (r_counter == (2047)) |
					      /**/
					      (r_counter == (2050)) |
					      /**/
					      (r_counter == (2053)) |
					      /**/
					      (r_counter == (2056)) |
					      /**/
					      (r_counter == (2059)) |
					      /**/
					      (r_counter == (2062)) |
					      /**/
					      (r_counter == (2065)) |
					      /**/
					      (r_counter == (2068)) |
					      /**/
					      (r_counter == (2071)) |
					      /**/
					      (r_counter == (2074)) |
					      /**/
					      (r_counter == (2077)) |
					      /**/
					      (r_counter == (2080)) |
					      /**/
					      (r_counter == (2083)) |
					      /**/
					      (r_counter == (2086)) |
					      /**/
					      (r_counter == (2089)) |
					      /**/
					      (r_counter == (2092)) |
					      /**/
					      (r_counter == (2095)) |
					      /**/
					      (r_counter == (2098)) |
					      /**/
					      (r_counter == (2101)) |
					      /**/
					      (r_counter == (2104)) |
					      /**/
					      (r_counter == (2107)) |
					      /**/
					      (r_counter == (2110)) |
					      /**/
					      (r_counter == (2113)) |
					      /**/
					      (r_counter == (2116)) |
					      /**/
					      (r_counter == (2119)) |
					      /**/
					      (r_counter == (2122)) |
					      /**/
					      (r_counter == (2125)) |
					      /**/
					      (r_counter == (2128)) |
					      /**/
					      (r_counter == (2131)) |
					      /**/
					      (r_counter == (2134)) |
					      /**/
					      (r_counter == (2137)) |
					      /**/
					      (r_counter == (2140)) |
					      /**/
					      (r_counter == (2143)) |
					      /**/
					      (r_counter == (2146)) |
					      /**/
					      (r_counter == (2149)) |
					      /**/
					      (r_counter == (2152)) |
					      /**/
					      (r_counter == (2155)) |
					      /**/
					      (r_counter == (2158)) |
					      /**/
					      (r_counter == (2161)) |
					      /**/
					      (r_counter == (2164)) |
					      /**/
					      (r_counter == (2167)) |
					      /**/
					      (r_counter == (2170)) |
					      /**/
					      (r_counter == (2173)) |
					      /**/
					      (r_counter == (2176)) |
					      /**/
					      (r_counter == (2179)) |
					      /**/
					      (r_counter == (2182)) |
					      /**/
					      (r_counter == (2185)) |
					      /**/
					      (r_counter == (2188)) |
					      /**/
					      (r_counter == (2191)) |
					      /**/
					      (r_counter == (2194)) |
					      /**/
					      (r_counter == (2197)) |
					      /**/
					      (r_counter == (2200)) |
					      /**/
					      (r_counter == (2203)) |
					      /**/
					      (r_counter == (2206)) |
					      /**/
					      (r_counter == (2209)) |
					      /**/
					      (r_counter == (2212)) |
					      /**/
					      (r_counter == (2215)) |
					      /**/
					      (r_counter == (2218)) |
					      /**/
					      (r_counter == (2221)) |
					      /**/
					      (r_counter == (2224)) |
					      /**/
					      (r_counter == (2227)) |
					      /**/
					      (r_counter == (2230)) |
					      /**/
					      (r_counter == (2233)) |
					      /**/
					      (r_counter == (2236)) |
					      /**/
					      (r_counter == (2239)) |
					      /**/
					      (r_counter == (2242)) |
					      /**/
					      (r_counter == (2245)) |
					      /**/
					      (r_counter == (2248)) |
					      /**/
					      (r_counter == (2251)) |
					      /**/
					      (r_counter == (2254)) |
					      /**/
					      (r_counter == (2257)) |
					      /**/
					      (r_counter == (2260)) |
					      /**/
					      (r_counter == (2263)) |
					      /**/
					      (r_counter == (2266)) |
					      /**/
					      (r_counter == (2269)) |
					      /**/
					      (r_counter == (2272)) |
					      /**/
					      (r_counter == (2275)) |
					      /**/
					      (r_counter == (2278)) |
					      /**/
					      (r_counter == (2281)) |
					      /**/
					      (r_counter == (2284)) |
					      /**/
					      (r_counter == (2287)) |
					      /**/
					      (r_counter == (2290)) |
					      /**/
					      (r_counter == (2293)) |
					      /**/
					      (r_counter == (2296)) |
					      /**/
					      (r_counter == (2299)) |
					      /**/
					      (r_counter == (2302)) |
					      /**/
					      (r_counter == (2305)) |
					      /**/
					      (r_counter == (2308)) |
					      /**/
					      (r_counter == (2311)) |
					      /**/
					      (r_counter == (2314)) |
					      /**/
					      (r_counter == (2317)) |
					      /**/
					      (r_counter == (2320)) |
					      /**/
					      (r_counter == (2323)) |
					      /**/
					      (r_counter == (2326)) |
					      /**/
					      (r_counter == (2329)) |
					      /**/
					      (r_counter == (2332)) |
					      /**/
					      (r_counter == (2335)) |
					      /**/
					      (r_counter == (2338)) |
					      /**/
					      (r_counter == (2341)) |
					      /**/
					      (r_counter == (2344)) |
					      /**/
					      (r_counter == (2347)) |
					      /**/
					      (r_counter == (2350)) |
					      /**/
					      (r_counter == (2353)) |
					      /**/
					      (r_counter == (2356)) |
					      /**/
					      (r_counter == (2359)) |
					      /**/
					      (r_counter == (2362)) |
					      /**/
					      (r_counter == (2365)) |
					      /**/
					      (r_counter == (2368)) |
					      /**/
					      (r_counter == (2371)) |
					      /**/
					      (r_counter == (2374)) |
					      /**/
					      (r_counter == (2377)) |
					      /**/
					      (r_counter == (2380)) |
					      /**/
					      (r_counter == (2383)) |
					      /**/
					      (r_counter == (2386)) |
					      /**/
					      (r_counter == (2389)) |
					      /**/
					      (r_counter == (2392)) |
					      /**/
					      (r_counter == (2395)) |
					      /**/
					      (r_counter == (2398)) |
					      /**/
					      (r_counter == (2401)));
   assign i_waddr_alpha=
			/**/
			(r_counter == (4)) ? 0:
			/**/
			(r_counter == (7)) ? 1:
			/**/
			(r_counter == (10)) ? 2:
			/**/
			(r_counter == (13)) ? 3:
			/**/
			(r_counter == (16)) ? 4:
			/**/
			(r_counter == (19)) ? 5:
			/**/
			(r_counter == (22)) ? 6:
			/**/
			(r_counter == (25)) ? 7:
			/**/
			(r_counter == (28)) ? 8:
			/**/
			(r_counter == (31)) ? 9:
			/**/
			(r_counter == (34)) ? 10:
			/**/
			(r_counter == (37)) ? 11:
			/**/
			(r_counter == (40)) ? 12:
			/**/
			(r_counter == (43)) ? 13:
			/**/
			(r_counter == (46)) ? 14:
			/**/
			(r_counter == (49)) ? 15:
			/**/
			(r_counter == (52)) ? 16:
			/**/
			(r_counter == (55)) ? 17:
			/**/
			(r_counter == (58)) ? 18:
			/**/
			(r_counter == (61)) ? 19:
			/**/
			(r_counter == (64)) ? 20:
			/**/
			(r_counter == (67)) ? 21:
			/**/
			(r_counter == (70)) ? 22:
			/**/
			(r_counter == (73)) ? 23:
			/**/
			(r_counter == (76)) ? 24:
			/**/
			(r_counter == (79)) ? 25:
			/**/
			(r_counter == (82)) ? 26:
			/**/
			(r_counter == (85)) ? 27:
			/**/
			(r_counter == (88)) ? 28:
			/**/
			(r_counter == (91)) ? 29:
			/**/
			(r_counter == (94)) ? 30:
			/**/
			(r_counter == (97)) ? 31:
			/**/
			(r_counter == (100)) ? 32:
			/**/
			(r_counter == (103)) ? 33:
			/**/
			(r_counter == (106)) ? 34:
			/**/
			(r_counter == (109)) ? 35:
			/**/
			(r_counter == (112)) ? 36:
			/**/
			(r_counter == (115)) ? 37:
			/**/
			(r_counter == (118)) ? 38:
			/**/
			(r_counter == (121)) ? 39:
			/**/
			(r_counter == (124)) ? 40:
			/**/
			(r_counter == (127)) ? 41:
			/**/
			(r_counter == (130)) ? 42:
			/**/
			(r_counter == (133)) ? 43:
			/**/
			(r_counter == (136)) ? 44:
			/**/
			(r_counter == (139)) ? 45:
			/**/
			(r_counter == (142)) ? 46:
			/**/
			(r_counter == (145)) ? 47:
			/**/
			(r_counter == (148)) ? 48:
			/**/
			(r_counter == (151)) ? 49:
			/**/
			(r_counter == (154)) ? 50:
			/**/
			(r_counter == (157)) ? 51:
			/**/
			(r_counter == (160)) ? 52:
			/**/
			(r_counter == (163)) ? 53:
			/**/
			(r_counter == (166)) ? 54:
			/**/
			(r_counter == (169)) ? 55:
			/**/
			(r_counter == (172)) ? 56:
			/**/
			(r_counter == (175)) ? 57:
			/**/
			(r_counter == (178)) ? 58:
			/**/
			(r_counter == (181)) ? 59:
			/**/
			(r_counter == (184)) ? 60:
			/**/
			(r_counter == (187)) ? 61:
			/**/
			(r_counter == (190)) ? 62:
			/**/
			(r_counter == (193)) ? 63:
			/**/
			(r_counter == (196)) ? 64:
			/**/
			(r_counter == (199)) ? 65:
			/**/
			(r_counter == (202)) ? 66:
			/**/
			(r_counter == (205)) ? 67:
			/**/
			(r_counter == (208)) ? 68:
			/**/
			(r_counter == (211)) ? 69:
			/**/
			(r_counter == (214)) ? 70:
			/**/
			(r_counter == (217)) ? 71:
			/**/
			(r_counter == (220)) ? 72:
			/**/
			(r_counter == (223)) ? 73:
			/**/
			(r_counter == (226)) ? 74:
			/**/
			(r_counter == (229)) ? 75:
			/**/
			(r_counter == (232)) ? 76:
			/**/
			(r_counter == (235)) ? 77:
			/**/
			(r_counter == (238)) ? 78:
			/**/
			(r_counter == (241)) ? 79:
			/**/
			(r_counter == (244)) ? 80:
			/**/
			(r_counter == (247)) ? 81:
			/**/
			(r_counter == (250)) ? 82:
			/**/
			(r_counter == (253)) ? 83:
			/**/
			(r_counter == (256)) ? 84:
			/**/
			(r_counter == (259)) ? 85:
			/**/
			(r_counter == (262)) ? 86:
			/**/
			(r_counter == (265)) ? 87:
			/**/
			(r_counter == (268)) ? 88:
			/**/
			(r_counter == (271)) ? 89:
			/**/
			(r_counter == (274)) ? 90:
			/**/
			(r_counter == (277)) ? 91:
			/**/
			(r_counter == (280)) ? 92:
			/**/
			(r_counter == (283)) ? 93:
			/**/
			(r_counter == (286)) ? 94:
			/**/
			(r_counter == (289)) ? 95:
			/**/
			(r_counter == (292)) ? 96:
			/**/
			(r_counter == (295)) ? 97:
			/**/
			(r_counter == (298)) ? 98:
			/**/
			(r_counter == (301)) ? 99:
			/**/
			(r_counter == (304)) ? 100:
			/**/
			(r_counter == (307)) ? 101:
			/**/
			(r_counter == (310)) ? 102:
			/**/
			(r_counter == (313)) ? 103:
			/**/
			(r_counter == (316)) ? 104:
			/**/
			(r_counter == (319)) ? 105:
			/**/
			(r_counter == (322)) ? 106:
			/**/
			(r_counter == (325)) ? 107:
			/**/
			(r_counter == (328)) ? 108:
			/**/
			(r_counter == (331)) ? 109:
			/**/
			(r_counter == (334)) ? 110:
			/**/
			(r_counter == (337)) ? 111:
			/**/
			(r_counter == (340)) ? 112:
			/**/
			(r_counter == (343)) ? 113:
			/**/
			(r_counter == (346)) ? 114:
			/**/
			(r_counter == (349)) ? 115:
			/**/
			(r_counter == (352)) ? 116:
			/**/
			(r_counter == (355)) ? 117:
			/**/
			(r_counter == (358)) ? 118:
			/**/
			(r_counter == (361)) ? 119:
			/**/
			(r_counter == (364)) ? 120:
			/**/
			(r_counter == (367)) ? 121:
			/**/
			(r_counter == (370)) ? 122:
			/**/
			(r_counter == (373)) ? 123:
			/**/
			(r_counter == (376)) ? 124:
			/**/
			(r_counter == (379)) ? 125:
			/**/
			(r_counter == (382)) ? 126:
			/**/
			(r_counter == (385)) ? 127:
			/**/
			(r_counter == (388)) ? 128:
			/**/
			(r_counter == (391)) ? 129:
			/**/
			(r_counter == (394)) ? 130:
			/**/
			(r_counter == (397)) ? 131:
			/**/
			(r_counter == (400)) ? 132:
			/**/
			(r_counter == (403)) ? 133:
			/**/
			(r_counter == (406)) ? 134:
			/**/
			(r_counter == (409)) ? 135:
			/**/
			(r_counter == (412)) ? 136:
			/**/
			(r_counter == (415)) ? 137:
			/**/
			(r_counter == (418)) ? 138:
			/**/
			(r_counter == (421)) ? 139:
			/**/
			(r_counter == (424)) ? 140:
			/**/
			(r_counter == (427)) ? 141:
			/**/
			(r_counter == (430)) ? 142:
			/**/
			(r_counter == (433)) ? 143:
			/**/
			(r_counter == (436)) ? 144:
			/**/
			(r_counter == (439)) ? 145:
			/**/
			(r_counter == (442)) ? 146:
			/**/
			(r_counter == (445)) ? 147:
			/**/
			(r_counter == (448)) ? 148:
			/**/
			(r_counter == (451)) ? 149:
			/**/
			(r_counter == (454)) ? 150:
			/**/
			(r_counter == (457)) ? 151:
			/**/
			(r_counter == (460)) ? 152:
			/**/
			(r_counter == (463)) ? 153:
			/**/
			(r_counter == (466)) ? 154:
			/**/
			(r_counter == (469)) ? 155:
			/**/
			(r_counter == (472)) ? 156:
			/**/
			(r_counter == (475)) ? 157:
			/**/
			(r_counter == (478)) ? 158:
			/**/
			(r_counter == (481)) ? 159:
			/**/
			(r_counter == (484)) ? 160:
			/**/
			(r_counter == (487)) ? 161:
			/**/
			(r_counter == (490)) ? 162:
			/**/
			(r_counter == (493)) ? 163:
			/**/
			(r_counter == (496)) ? 164:
			/**/
			(r_counter == (499)) ? 165:
			/**/
			(r_counter == (502)) ? 166:
			/**/
			(r_counter == (505)) ? 167:
			/**/
			(r_counter == (508)) ? 168:
			/**/
			(r_counter == (511)) ? 169:
			/**/
			(r_counter == (514)) ? 170:
			/**/
			(r_counter == (517)) ? 171:
			/**/
			(r_counter == (520)) ? 172:
			/**/
			(r_counter == (523)) ? 173:
			/**/
			(r_counter == (526)) ? 174:
			/**/
			(r_counter == (529)) ? 175:
			/**/
			(r_counter == (532)) ? 176:
			/**/
			(r_counter == (535)) ? 177:
			/**/
			(r_counter == (538)) ? 178:
			/**/
			(r_counter == (541)) ? 179:
			/**/
			(r_counter == (544)) ? 180:
			/**/
			(r_counter == (547)) ? 181:
			/**/
			(r_counter == (550)) ? 182:
			/**/
			(r_counter == (553)) ? 183:
			/**/
			(r_counter == (556)) ? 184:
			/**/
			(r_counter == (559)) ? 185:
			/**/
			(r_counter == (562)) ? 186:
			/**/
			(r_counter == (565)) ? 187:
			/**/
			(r_counter == (568)) ? 188:
			/**/
			(r_counter == (571)) ? 189:
			/**/
			(r_counter == (574)) ? 190:
			/**/
			(r_counter == (577)) ? 191:
			/**/
			(r_counter == (580)) ? 192:
			/**/
			(r_counter == (583)) ? 193:
			/**/
			(r_counter == (586)) ? 194:
			/**/
			(r_counter == (589)) ? 195:
			/**/
			(r_counter == (592)) ? 196:
			/**/
			(r_counter == (595)) ? 197:
			/**/
			(r_counter == (598)) ? 198:
			/**/
			(r_counter == (601)) ? 199:
			/**/
			(r_counter == (604)) ? 200:
			/**/
			(r_counter == (607)) ? 201:
			/**/
			(r_counter == (610)) ? 202:
			/**/
			(r_counter == (613)) ? 203:
			/**/
			(r_counter == (616)) ? 204:
			/**/
			(r_counter == (619)) ? 205:
			/**/
			(r_counter == (622)) ? 206:
			/**/
			(r_counter == (625)) ? 207:
			/**/
			(r_counter == (628)) ? 208:
			/**/
			(r_counter == (631)) ? 209:
			/**/
			(r_counter == (634)) ? 210:
			/**/
			(r_counter == (637)) ? 211:
			/**/
			(r_counter == (640)) ? 212:
			/**/
			(r_counter == (643)) ? 213:
			/**/
			(r_counter == (646)) ? 214:
			/**/
			(r_counter == (649)) ? 215:
			/**/
			(r_counter == (652)) ? 216:
			/**/
			(r_counter == (655)) ? 217:
			/**/
			(r_counter == (658)) ? 218:
			/**/
			(r_counter == (661)) ? 219:
			/**/
			(r_counter == (664)) ? 220:
			/**/
			(r_counter == (667)) ? 221:
			/**/
			(r_counter == (670)) ? 222:
			/**/
			(r_counter == (673)) ? 223:
			/**/
			(r_counter == (676)) ? 224:
			/**/
			(r_counter == (679)) ? 225:
			/**/
			(r_counter == (682)) ? 226:
			/**/
			(r_counter == (685)) ? 227:
			/**/
			(r_counter == (688)) ? 228:
			/**/
			(r_counter == (691)) ? 229:
			/**/
			(r_counter == (694)) ? 230:
			/**/
			(r_counter == (697)) ? 231:
			/**/
			(r_counter == (700)) ? 232:
			/**/
			(r_counter == (703)) ? 233:
			/**/
			(r_counter == (706)) ? 234:
			/**/
			(r_counter == (709)) ? 235:
			/**/
			(r_counter == (712)) ? 236:
			/**/
			(r_counter == (715)) ? 237:
			/**/
			(r_counter == (718)) ? 238:
			/**/
			(r_counter == (721)) ? 239:
			/**/
			(r_counter == (724)) ? 240:
			/**/
			(r_counter == (727)) ? 241:
			/**/
			(r_counter == (730)) ? 242:
			/**/
			(r_counter == (733)) ? 243:
			/**/
			(r_counter == (736)) ? 244:
			/**/
			(r_counter == (739)) ? 245:
			/**/
			(r_counter == (742)) ? 246:
			/**/
			(r_counter == (745)) ? 247:
			/**/
			(r_counter == (748)) ? 248:
			/**/
			(r_counter == (751)) ? 249:
			/**/
			(r_counter == (754)) ? 250:
			/**/
			(r_counter == (757)) ? 251:
			/**/
			(r_counter == (760)) ? 252:
			/**/
			(r_counter == (763)) ? 253:
			/**/
			(r_counter == (766)) ? 254:
			/**/
			(r_counter == (769)) ? 255:
			/**/
			(r_counter == (772)) ? 256:
			/**/
			(r_counter == (775)) ? 257:
			/**/
			(r_counter == (778)) ? 258:
			/**/
			(r_counter == (781)) ? 259:
			/**/
			(r_counter == (784)) ? 260:
			/**/
			(r_counter == (787)) ? 261:
			/**/
			(r_counter == (790)) ? 262:
			/**/
			(r_counter == (793)) ? 263:
			/**/
			(r_counter == (796)) ? 264:
			/**/
			(r_counter == (799)) ? 265:
			/**/
			(r_counter == (802)) ? 266:
			/**/
			(r_counter == (805)) ? 267:
			/**/
			(r_counter == (808)) ? 268:
			/**/
			(r_counter == (811)) ? 269:
			/**/
			(r_counter == (814)) ? 270:
			/**/
			(r_counter == (817)) ? 271:
			/**/
			(r_counter == (820)) ? 272:
			/**/
			(r_counter == (823)) ? 273:
			/**/
			(r_counter == (826)) ? 274:
			/**/
			(r_counter == (829)) ? 275:
			/**/
			(r_counter == (832)) ? 276:
			/**/
			(r_counter == (835)) ? 277:
			/**/
			(r_counter == (838)) ? 278:
			/**/
			(r_counter == (841)) ? 279:
			/**/
			(r_counter == (844)) ? 280:
			/**/
			(r_counter == (847)) ? 281:
			/**/
			(r_counter == (850)) ? 282:
			/**/
			(r_counter == (853)) ? 283:
			/**/
			(r_counter == (856)) ? 284:
			/**/
			(r_counter == (859)) ? 285:
			/**/
			(r_counter == (862)) ? 286:
			/**/
			(r_counter == (865)) ? 287:
			/**/
			(r_counter == (868)) ? 288:
			/**/
			(r_counter == (871)) ? 289:
			/**/
			(r_counter == (874)) ? 290:
			/**/
			(r_counter == (877)) ? 291:
			/**/
			(r_counter == (880)) ? 292:
			/**/
			(r_counter == (883)) ? 293:
			/**/
			(r_counter == (886)) ? 294:
			/**/
			(r_counter == (889)) ? 295:
			/**/
			(r_counter == (892)) ? 296:
			/**/
			(r_counter == (895)) ? 297:
			/**/
			(r_counter == (898)) ? 298:
			/**/
			(r_counter == (901)) ? 299:
			/**/
			(r_counter == (904)) ? 300:
			/**/
			(r_counter == (907)) ? 301:
			/**/
			(r_counter == (910)) ? 302:
			/**/
			(r_counter == (913)) ? 303:
			/**/
			(r_counter == (916)) ? 304:
			/**/
			(r_counter == (919)) ? 305:
			/**/
			(r_counter == (922)) ? 306:
			/**/
			(r_counter == (925)) ? 307:
			/**/
			(r_counter == (928)) ? 308:
			/**/
			(r_counter == (931)) ? 309:
			/**/
			(r_counter == (934)) ? 310:
			/**/
			(r_counter == (937)) ? 311:
			/**/
			(r_counter == (940)) ? 312:
			/**/
			(r_counter == (943)) ? 313:
			/**/
			(r_counter == (946)) ? 314:
			/**/
			(r_counter == (949)) ? 315:
			/**/
			(r_counter == (952)) ? 316:
			/**/
			(r_counter == (955)) ? 317:
			/**/
			(r_counter == (958)) ? 318:
			/**/
			(r_counter == (961)) ? 319:
			/**/
			(r_counter == (964)) ? 320:
			/**/
			(r_counter == (967)) ? 321:
			/**/
			(r_counter == (970)) ? 322:
			/**/
			(r_counter == (973)) ? 323:
			/**/
			(r_counter == (976)) ? 324:
			/**/
			(r_counter == (979)) ? 325:
			/**/
			(r_counter == (982)) ? 326:
			/**/
			(r_counter == (985)) ? 327:
			/**/
			(r_counter == (988)) ? 328:
			/**/
			(r_counter == (991)) ? 329:
			/**/
			(r_counter == (994)) ? 330:
			/**/
			(r_counter == (997)) ? 331:
			/**/
			(r_counter == (1000)) ? 332:
			/**/
			(r_counter == (1003)) ? 333:
			/**/
			(r_counter == (1006)) ? 334:
			/**/
			(r_counter == (1009)) ? 335:
			/**/
			(r_counter == (1012)) ? 336:
			/**/
			(r_counter == (1015)) ? 337:
			/**/
			(r_counter == (1018)) ? 338:
			/**/
			(r_counter == (1021)) ? 339:
			/**/
			(r_counter == (1024)) ? 340:
			/**/
			(r_counter == (1027)) ? 341:
			/**/
			(r_counter == (1030)) ? 342:
			/**/
			(r_counter == (1033)) ? 343:
			/**/
			(r_counter == (1036)) ? 344:
			/**/
			(r_counter == (1039)) ? 345:
			/**/
			(r_counter == (1042)) ? 346:
			/**/
			(r_counter == (1045)) ? 347:
			/**/
			(r_counter == (1048)) ? 348:
			/**/
			(r_counter == (1051)) ? 349:
			/**/
			(r_counter == (1054)) ? 350:
			/**/
			(r_counter == (1057)) ? 351:
			/**/
			(r_counter == (1060)) ? 352:
			/**/
			(r_counter == (1063)) ? 353:
			/**/
			(r_counter == (1066)) ? 354:
			/**/
			(r_counter == (1069)) ? 355:
			/**/
			(r_counter == (1072)) ? 356:
			/**/
			(r_counter == (1075)) ? 357:
			/**/
			(r_counter == (1078)) ? 358:
			/**/
			(r_counter == (1081)) ? 359:
			/**/
			(r_counter == (1084)) ? 360:
			/**/
			(r_counter == (1087)) ? 361:
			/**/
			(r_counter == (1090)) ? 362:
			/**/
			(r_counter == (1093)) ? 363:
			/**/
			(r_counter == (1096)) ? 364:
			/**/
			(r_counter == (1099)) ? 365:
			/**/
			(r_counter == (1102)) ? 366:
			/**/
			(r_counter == (1105)) ? 367:
			/**/
			(r_counter == (1108)) ? 368:
			/**/
			(r_counter == (1111)) ? 369:
			/**/
			(r_counter == (1114)) ? 370:
			/**/
			(r_counter == (1117)) ? 371:
			/**/
			(r_counter == (1120)) ? 372:
			/**/
			(r_counter == (1123)) ? 373:
			/**/
			(r_counter == (1126)) ? 374:
			/**/
			(r_counter == (1129)) ? 375:
			/**/
			(r_counter == (1132)) ? 376:
			/**/
			(r_counter == (1135)) ? 377:
			/**/
			(r_counter == (1138)) ? 378:
			/**/
			(r_counter == (1141)) ? 379:
			/**/
			(r_counter == (1144)) ? 380:
			/**/
			(r_counter == (1147)) ? 381:
			/**/
			(r_counter == (1150)) ? 382:
			/**/
			(r_counter == (1153)) ? 383:
			/**/
			(r_counter == (1156)) ? 384:
			/**/
			(r_counter == (1159)) ? 385:
			/**/
			(r_counter == (1162)) ? 386:
			/**/
			(r_counter == (1165)) ? 387:
			/**/
			(r_counter == (1168)) ? 388:
			/**/
			(r_counter == (1171)) ? 389:
			/**/
			(r_counter == (1174)) ? 390:
			/**/
			(r_counter == (1177)) ? 391:
			/**/
			(r_counter == (1180)) ? 392:
			/**/
			(r_counter == (1183)) ? 393:
			/**/
			(r_counter == (1186)) ? 394:
			/**/
			(r_counter == (1189)) ? 395:
			/**/
			(r_counter == (1192)) ? 396:
			/**/
			(r_counter == (1195)) ? 397:
			/**/
			(r_counter == (1198)) ? 398:
			/**/
			(r_counter == (1201)) ? 399:
			/**/
			(r_counter == (1204)) ? 400:
			/**/
			(r_counter == (1207)) ? 401:
			/**/
			(r_counter == (1210)) ? 402:
			/**/
			(r_counter == (1213)) ? 403:
			/**/
			(r_counter == (1216)) ? 404:
			/**/
			(r_counter == (1219)) ? 405:
			/**/
			(r_counter == (1222)) ? 406:
			/**/
			(r_counter == (1225)) ? 407:
			/**/
			(r_counter == (1228)) ? 408:
			/**/
			(r_counter == (1231)) ? 409:
			/**/
			(r_counter == (1234)) ? 410:
			/**/
			(r_counter == (1237)) ? 411:
			/**/
			(r_counter == (1240)) ? 412:
			/**/
			(r_counter == (1243)) ? 413:
			/**/
			(r_counter == (1246)) ? 414:
			/**/
			(r_counter == (1249)) ? 415:
			/**/
			(r_counter == (1252)) ? 416:
			/**/
			(r_counter == (1255)) ? 417:
			/**/
			(r_counter == (1258)) ? 418:
			/**/
			(r_counter == (1261)) ? 419:
			/**/
			(r_counter == (1264)) ? 420:
			/**/
			(r_counter == (1267)) ? 421:
			/**/
			(r_counter == (1270)) ? 422:
			/**/
			(r_counter == (1273)) ? 423:
			/**/
			(r_counter == (1276)) ? 424:
			/**/
			(r_counter == (1279)) ? 425:
			/**/
			(r_counter == (1282)) ? 426:
			/**/
			(r_counter == (1285)) ? 427:
			/**/
			(r_counter == (1288)) ? 428:
			/**/
			(r_counter == (1291)) ? 429:
			/**/
			(r_counter == (1294)) ? 430:
			/**/
			(r_counter == (1297)) ? 431:
			/**/
			(r_counter == (1300)) ? 432:
			/**/
			(r_counter == (1303)) ? 433:
			/**/
			(r_counter == (1306)) ? 434:
			/**/
			(r_counter == (1309)) ? 435:
			/**/
			(r_counter == (1312)) ? 436:
			/**/
			(r_counter == (1315)) ? 437:
			/**/
			(r_counter == (1318)) ? 438:
			/**/
			(r_counter == (1321)) ? 439:
			/**/
			(r_counter == (1324)) ? 440:
			/**/
			(r_counter == (1327)) ? 441:
			/**/
			(r_counter == (1330)) ? 442:
			/**/
			(r_counter == (1333)) ? 443:
			/**/
			(r_counter == (1336)) ? 444:
			/**/
			(r_counter == (1339)) ? 445:
			/**/
			(r_counter == (1342)) ? 446:
			/**/
			(r_counter == (1345)) ? 447:
			/**/
			(r_counter == (1348)) ? 448:
			/**/
			(r_counter == (1351)) ? 449:
			/**/
			(r_counter == (1354)) ? 450:
			/**/
			(r_counter == (1357)) ? 451:
			/**/
			(r_counter == (1360)) ? 452:
			/**/
			(r_counter == (1363)) ? 453:
			/**/
			(r_counter == (1366)) ? 454:
			/**/
			(r_counter == (1369)) ? 455:
			/**/
			(r_counter == (1372)) ? 456:
			/**/
			(r_counter == (1375)) ? 457:
			/**/
			(r_counter == (1378)) ? 458:
			/**/
			(r_counter == (1381)) ? 459:
			/**/
			(r_counter == (1384)) ? 460:
			/**/
			(r_counter == (1387)) ? 461:
			/**/
			(r_counter == (1390)) ? 462:
			/**/
			(r_counter == (1393)) ? 463:
			/**/
			(r_counter == (1396)) ? 464:
			/**/
			(r_counter == (1399)) ? 465:
			/**/
			(r_counter == (1402)) ? 466:
			/**/
			(r_counter == (1405)) ? 467:
			/**/
			(r_counter == (1408)) ? 468:
			/**/
			(r_counter == (1411)) ? 469:
			/**/
			(r_counter == (1414)) ? 470:
			/**/
			(r_counter == (1417)) ? 471:
			/**/
			(r_counter == (1420)) ? 472:
			/**/
			(r_counter == (1423)) ? 473:
			/**/
			(r_counter == (1426)) ? 474:
			/**/
			(r_counter == (1429)) ? 475:
			/**/
			(r_counter == (1432)) ? 476:
			/**/
			(r_counter == (1435)) ? 477:
			/**/
			(r_counter == (1438)) ? 478:
			/**/
			(r_counter == (1441)) ? 479:
			/**/
			(r_counter == (1444)) ? 480:
			/**/
			(r_counter == (1447)) ? 481:
			/**/
			(r_counter == (1450)) ? 482:
			/**/
			(r_counter == (1453)) ? 483:
			/**/
			(r_counter == (1456)) ? 484:
			/**/
			(r_counter == (1459)) ? 485:
			/**/
			(r_counter == (1462)) ? 486:
			/**/
			(r_counter == (1465)) ? 487:
			/**/
			(r_counter == (1468)) ? 488:
			/**/
			(r_counter == (1471)) ? 489:
			/**/
			(r_counter == (1474)) ? 490:
			/**/
			(r_counter == (1477)) ? 491:
			/**/
			(r_counter == (1480)) ? 492:
			/**/
			(r_counter == (1483)) ? 493:
			/**/
			(r_counter == (1486)) ? 494:
			/**/
			(r_counter == (1489)) ? 495:
			/**/
			(r_counter == (1492)) ? 496:
			/**/
			(r_counter == (1495)) ? 497:
			/**/
			(r_counter == (1498)) ? 498:
			/**/
			(r_counter == (1501)) ? 499:
			/**/
			(r_counter == (1504)) ? 500:
			/**/
			(r_counter == (1507)) ? 501:
			/**/
			(r_counter == (1510)) ? 502:
			/**/
			(r_counter == (1513)) ? 503:
			/**/
			(r_counter == (1516)) ? 504:
			/**/
			(r_counter == (1519)) ? 505:
			/**/
			(r_counter == (1522)) ? 506:
			/**/
			(r_counter == (1525)) ? 507:
			/**/
			(r_counter == (1528)) ? 508:
			/**/
			(r_counter == (1531)) ? 509:
			/**/
			(r_counter == (1534)) ? 510:
			/**/
			(r_counter == (1537)) ? 511:
			/**/
			(r_counter == (1540)) ? 512:
			/**/
			(r_counter == (1543)) ? 513:
			/**/
			(r_counter == (1546)) ? 514:
			/**/
			(r_counter == (1549)) ? 515:
			/**/
			(r_counter == (1552)) ? 516:
			/**/
			(r_counter == (1555)) ? 517:
			/**/
			(r_counter == (1558)) ? 518:
			/**/
			(r_counter == (1561)) ? 519:
			/**/
			(r_counter == (1564)) ? 520:
			/**/
			(r_counter == (1567)) ? 521:
			/**/
			(r_counter == (1570)) ? 522:
			/**/
			(r_counter == (1573)) ? 523:
			/**/
			(r_counter == (1576)) ? 524:
			/**/
			(r_counter == (1579)) ? 525:
			/**/
			(r_counter == (1582)) ? 526:
			/**/
			(r_counter == (1585)) ? 527:
			/**/
			(r_counter == (1588)) ? 528:
			/**/
			(r_counter == (1591)) ? 529:
			/**/
			(r_counter == (1594)) ? 530:
			/**/
			(r_counter == (1597)) ? 531:
			/**/
			(r_counter == (1600)) ? 532:
			/**/
			(r_counter == (1603)) ? 533:
			/**/
			(r_counter == (1606)) ? 534:
			/**/
			(r_counter == (1609)) ? 535:
			/**/
			(r_counter == (1612)) ? 536:
			/**/
			(r_counter == (1615)) ? 537:
			/**/
			(r_counter == (1618)) ? 538:
			/**/
			(r_counter == (1621)) ? 539:
			/**/
			(r_counter == (1624)) ? 540:
			/**/
			(r_counter == (1627)) ? 541:
			/**/
			(r_counter == (1630)) ? 542:
			/**/
			(r_counter == (1633)) ? 543:
			/**/
			(r_counter == (1636)) ? 544:
			/**/
			(r_counter == (1639)) ? 545:
			/**/
			(r_counter == (1642)) ? 546:
			/**/
			(r_counter == (1645)) ? 547:
			/**/
			(r_counter == (1648)) ? 548:
			/**/
			(r_counter == (1651)) ? 549:
			/**/
			(r_counter == (1654)) ? 550:
			/**/
			(r_counter == (1657)) ? 551:
			/**/
			(r_counter == (1660)) ? 552:
			/**/
			(r_counter == (1663)) ? 553:
			/**/
			(r_counter == (1666)) ? 554:
			/**/
			(r_counter == (1669)) ? 555:
			/**/
			(r_counter == (1672)) ? 556:
			/**/
			(r_counter == (1675)) ? 557:
			/**/
			(r_counter == (1678)) ? 558:
			/**/
			(r_counter == (1681)) ? 559:
			/**/
			(r_counter == (1684)) ? 560:
			/**/
			(r_counter == (1687)) ? 561:
			/**/
			(r_counter == (1690)) ? 562:
			/**/
			(r_counter == (1693)) ? 563:
			/**/
			(r_counter == (1696)) ? 564:
			/**/
			(r_counter == (1699)) ? 565:
			/**/
			(r_counter == (1702)) ? 566:
			/**/
			(r_counter == (1705)) ? 567:
			/**/
			(r_counter == (1708)) ? 568:
			/**/
			(r_counter == (1711)) ? 569:
			/**/
			(r_counter == (1714)) ? 570:
			/**/
			(r_counter == (1717)) ? 571:
			/**/
			(r_counter == (1720)) ? 572:
			/**/
			(r_counter == (1723)) ? 573:
			/**/
			(r_counter == (1726)) ? 574:
			/**/
			(r_counter == (1729)) ? 575:
			/**/
			(r_counter == (1732)) ? 576:
			/**/
			(r_counter == (1735)) ? 577:
			/**/
			(r_counter == (1738)) ? 578:
			/**/
			(r_counter == (1741)) ? 579:
			/**/
			(r_counter == (1744)) ? 580:
			/**/
			(r_counter == (1747)) ? 581:
			/**/
			(r_counter == (1750)) ? 582:
			/**/
			(r_counter == (1753)) ? 583:
			/**/
			(r_counter == (1756)) ? 584:
			/**/
			(r_counter == (1759)) ? 585:
			/**/
			(r_counter == (1762)) ? 586:
			/**/
			(r_counter == (1765)) ? 587:
			/**/
			(r_counter == (1768)) ? 588:
			/**/
			(r_counter == (1771)) ? 589:
			/**/
			(r_counter == (1774)) ? 590:
			/**/
			(r_counter == (1777)) ? 591:
			/**/
			(r_counter == (1780)) ? 592:
			/**/
			(r_counter == (1783)) ? 593:
			/**/
			(r_counter == (1786)) ? 594:
			/**/
			(r_counter == (1789)) ? 595:
			/**/
			(r_counter == (1792)) ? 596:
			/**/
			(r_counter == (1795)) ? 597:
			/**/
			(r_counter == (1798)) ? 598:
			/**/
			(r_counter == (1801)) ? 599:
			/**/
			(r_counter == (1804)) ? 600:
			/**/
			(r_counter == (1807)) ? 601:
			/**/
			(r_counter == (1810)) ? 602:
			/**/
			(r_counter == (1813)) ? 603:
			/**/
			(r_counter == (1816)) ? 604:
			/**/
			(r_counter == (1819)) ? 605:
			/**/
			(r_counter == (1822)) ? 606:
			/**/
			(r_counter == (1825)) ? 607:
			/**/
			(r_counter == (1828)) ? 608:
			/**/
			(r_counter == (1831)) ? 609:
			/**/
			(r_counter == (1834)) ? 610:
			/**/
			(r_counter == (1837)) ? 611:
			/**/
			(r_counter == (1840)) ? 612:
			/**/
			(r_counter == (1843)) ? 613:
			/**/
			(r_counter == (1846)) ? 614:
			/**/
			(r_counter == (1849)) ? 615:
			/**/
			(r_counter == (1852)) ? 616:
			/**/
			(r_counter == (1855)) ? 617:
			/**/
			(r_counter == (1858)) ? 618:
			/**/
			(r_counter == (1861)) ? 619:
			/**/
			(r_counter == (1864)) ? 620:
			/**/
			(r_counter == (1867)) ? 621:
			/**/
			(r_counter == (1870)) ? 622:
			/**/
			(r_counter == (1873)) ? 623:
			/**/
			(r_counter == (1876)) ? 624:
			/**/
			(r_counter == (1879)) ? 625:
			/**/
			(r_counter == (1882)) ? 626:
			/**/
			(r_counter == (1885)) ? 627:
			/**/
			(r_counter == (1888)) ? 628:
			/**/
			(r_counter == (1891)) ? 629:
			/**/
			(r_counter == (1894)) ? 630:
			/**/
			(r_counter == (1897)) ? 631:
			/**/
			(r_counter == (1900)) ? 632:
			/**/
			(r_counter == (1903)) ? 633:
			/**/
			(r_counter == (1906)) ? 634:
			/**/
			(r_counter == (1909)) ? 635:
			/**/
			(r_counter == (1912)) ? 636:
			/**/
			(r_counter == (1915)) ? 637:
			/**/
			(r_counter == (1918)) ? 638:
			/**/
			(r_counter == (1921)) ? 639:
			/**/
			(r_counter == (1924)) ? 640:
			/**/
			(r_counter == (1927)) ? 641:
			/**/
			(r_counter == (1930)) ? 642:
			/**/
			(r_counter == (1933)) ? 643:
			/**/
			(r_counter == (1936)) ? 644:
			/**/
			(r_counter == (1939)) ? 645:
			/**/
			(r_counter == (1942)) ? 646:
			/**/
			(r_counter == (1945)) ? 647:
			/**/
			(r_counter == (1948)) ? 648:
			/**/
			(r_counter == (1951)) ? 649:
			/**/
			(r_counter == (1954)) ? 650:
			/**/
			(r_counter == (1957)) ? 651:
			/**/
			(r_counter == (1960)) ? 652:
			/**/
			(r_counter == (1963)) ? 653:
			/**/
			(r_counter == (1966)) ? 654:
			/**/
			(r_counter == (1969)) ? 655:
			/**/
			(r_counter == (1972)) ? 656:
			/**/
			(r_counter == (1975)) ? 657:
			/**/
			(r_counter == (1978)) ? 658:
			/**/
			(r_counter == (1981)) ? 659:
			/**/
			(r_counter == (1984)) ? 660:
			/**/
			(r_counter == (1987)) ? 661:
			/**/
			(r_counter == (1990)) ? 662:
			/**/
			(r_counter == (1993)) ? 663:
			/**/
			(r_counter == (1996)) ? 664:
			/**/
			(r_counter == (1999)) ? 665:
			/**/
			(r_counter == (2002)) ? 666:
			/**/
			(r_counter == (2005)) ? 667:
			/**/
			(r_counter == (2008)) ? 668:
			/**/
			(r_counter == (2011)) ? 669:
			/**/
			(r_counter == (2014)) ? 670:
			/**/
			(r_counter == (2017)) ? 671:
			/**/
			(r_counter == (2020)) ? 672:
			/**/
			(r_counter == (2023)) ? 673:
			/**/
			(r_counter == (2026)) ? 674:
			/**/
			(r_counter == (2029)) ? 675:
			/**/
			(r_counter == (2032)) ? 676:
			/**/
			(r_counter == (2035)) ? 677:
			/**/
			(r_counter == (2038)) ? 678:
			/**/
			(r_counter == (2041)) ? 679:
			/**/
			(r_counter == (2044)) ? 680:
			/**/
			(r_counter == (2047)) ? 681:
			/**/
			(r_counter == (2050)) ? 682:
			/**/
			(r_counter == (2053)) ? 683:
			/**/
			(r_counter == (2056)) ? 684:
			/**/
			(r_counter == (2059)) ? 685:
			/**/
			(r_counter == (2062)) ? 686:
			/**/
			(r_counter == (2065)) ? 687:
			/**/
			(r_counter == (2068)) ? 688:
			/**/
			(r_counter == (2071)) ? 689:
			/**/
			(r_counter == (2074)) ? 690:
			/**/
			(r_counter == (2077)) ? 691:
			/**/
			(r_counter == (2080)) ? 692:
			/**/
			(r_counter == (2083)) ? 693:
			/**/
			(r_counter == (2086)) ? 694:
			/**/
			(r_counter == (2089)) ? 695:
			/**/
			(r_counter == (2092)) ? 696:
			/**/
			(r_counter == (2095)) ? 697:
			/**/
			(r_counter == (2098)) ? 698:
			/**/
			(r_counter == (2101)) ? 699:
			/**/
			(r_counter == (2104)) ? 700:
			/**/
			(r_counter == (2107)) ? 701:
			/**/
			(r_counter == (2110)) ? 702:
			/**/
			(r_counter == (2113)) ? 703:
			/**/
			(r_counter == (2116)) ? 704:
			/**/
			(r_counter == (2119)) ? 705:
			/**/
			(r_counter == (2122)) ? 706:
			/**/
			(r_counter == (2125)) ? 707:
			/**/
			(r_counter == (2128)) ? 708:
			/**/
			(r_counter == (2131)) ? 709:
			/**/
			(r_counter == (2134)) ? 710:
			/**/
			(r_counter == (2137)) ? 711:
			/**/
			(r_counter == (2140)) ? 712:
			/**/
			(r_counter == (2143)) ? 713:
			/**/
			(r_counter == (2146)) ? 714:
			/**/
			(r_counter == (2149)) ? 715:
			/**/
			(r_counter == (2152)) ? 716:
			/**/
			(r_counter == (2155)) ? 717:
			/**/
			(r_counter == (2158)) ? 718:
			/**/
			(r_counter == (2161)) ? 719:
			/**/
			(r_counter == (2164)) ? 720:
			/**/
			(r_counter == (2167)) ? 721:
			/**/
			(r_counter == (2170)) ? 722:
			/**/
			(r_counter == (2173)) ? 723:
			/**/
			(r_counter == (2176)) ? 724:
			/**/
			(r_counter == (2179)) ? 725:
			/**/
			(r_counter == (2182)) ? 726:
			/**/
			(r_counter == (2185)) ? 727:
			/**/
			(r_counter == (2188)) ? 728:
			/**/
			(r_counter == (2191)) ? 729:
			/**/
			(r_counter == (2194)) ? 730:
			/**/
			(r_counter == (2197)) ? 731:
			/**/
			(r_counter == (2200)) ? 732:
			/**/
			(r_counter == (2203)) ? 733:
			/**/
			(r_counter == (2206)) ? 734:
			/**/
			(r_counter == (2209)) ? 735:
			/**/
			(r_counter == (2212)) ? 736:
			/**/
			(r_counter == (2215)) ? 737:
			/**/
			(r_counter == (2218)) ? 738:
			/**/
			(r_counter == (2221)) ? 739:
			/**/
			(r_counter == (2224)) ? 740:
			/**/
			(r_counter == (2227)) ? 741:
			/**/
			(r_counter == (2230)) ? 742:
			/**/
			(r_counter == (2233)) ? 743:
			/**/
			(r_counter == (2236)) ? 744:
			/**/
			(r_counter == (2239)) ? 745:
			/**/
			(r_counter == (2242)) ? 746:
			/**/
			(r_counter == (2245)) ? 747:
			/**/
			(r_counter == (2248)) ? 748:
			/**/
			(r_counter == (2251)) ? 749:
			/**/
			(r_counter == (2254)) ? 750:
			/**/
			(r_counter == (2257)) ? 751:
			/**/
			(r_counter == (2260)) ? 752:
			/**/
			(r_counter == (2263)) ? 753:
			/**/
			(r_counter == (2266)) ? 754:
			/**/
			(r_counter == (2269)) ? 755:
			/**/
			(r_counter == (2272)) ? 756:
			/**/
			(r_counter == (2275)) ? 757:
			/**/
			(r_counter == (2278)) ? 758:
			/**/
			(r_counter == (2281)) ? 759:
			/**/
			(r_counter == (2284)) ? 760:
			/**/
			(r_counter == (2287)) ? 761:
			/**/
			(r_counter == (2290)) ? 762:
			/**/
			(r_counter == (2293)) ? 763:
			/**/
			(r_counter == (2296)) ? 764:
			/**/
			(r_counter == (2299)) ? 765:
			/**/
			(r_counter == (2302)) ? 766:
			/**/
			(r_counter == (2305)) ? 767:
			/**/
			(r_counter == (2308)) ? 768:
			/**/
			(r_counter == (2311)) ? 769:
			/**/
			(r_counter == (2314)) ? 770:
			/**/
			(r_counter == (2317)) ? 771:
			/**/
			(r_counter == (2320)) ? 772:
			/**/
			(r_counter == (2323)) ? 773:
			/**/
			(r_counter == (2326)) ? 774:
			/**/
			(r_counter == (2329)) ? 775:
			/**/
			(r_counter == (2332)) ? 776:
			/**/
			(r_counter == (2335)) ? 777:
			/**/
			(r_counter == (2338)) ? 778:
			/**/
			(r_counter == (2341)) ? 779:
			/**/
			(r_counter == (2344)) ? 780:
			/**/
			(r_counter == (2347)) ? 781:
			/**/
			(r_counter == (2350)) ? 782:
			/**/
			(r_counter == (2353)) ? 783:
			/**/
			(r_counter == (2356)) ? 784:
			/**/
			(r_counter == (2359)) ? 785:
			/**/
			(r_counter == (2362)) ? 786:
			/**/
			(r_counter == (2365)) ? 787:
			/**/
			(r_counter == (2368)) ? 788:
			/**/
			(r_counter == (2371)) ? 789:
			/**/
			(r_counter == (2374)) ? 790:
			/**/
			(r_counter == (2377)) ? 791:
			/**/
			(r_counter == (2380)) ? 792:
			/**/
			(r_counter == (2383)) ? 793:
			/**/
			(r_counter == (2386)) ? 794:
			/**/
			(r_counter == (2389)) ? 795:
			/**/
			(r_counter == (2392)) ? 796:
			/**/
			(r_counter == (2395)) ? 797:
			/**/
			(r_counter == (2398)) ? 798:
			/**/
			(r_counter == (2401)) ? 799:
			/**/
			(r_counter == (2404)) ? 800:
			/**/
			0;
   
   assign i_raddr_alpha=/**/
		        /**/ 
			(r_counter == 0 & r_state==zStateColumn) ? 565:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 2 & r_state==zStateColumn) ? 566:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 4 & r_state==zStateColumn) ? 489:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 6 & r_state==zStateColumn) ? 678:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 8 & r_state==zStateColumn) ? 794:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 10 & r_state==zStateColumn) ? 404:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 12 & r_state==zStateColumn) ? 509:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 14 & r_state==zStateColumn) ? 422:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 16 & r_state==zStateColumn) ? 642:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 18 & r_state==zStateColumn) ? 561:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 20 & r_state==zStateColumn) ? 434:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 22 & r_state==zStateColumn) ? 657:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 24 & r_state==zStateColumn) ? 517:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 26 & r_state==zStateColumn) ? 537:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 28 & r_state==zStateColumn) ? 554:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 30 & r_state==zStateColumn) ? 766:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 32 & r_state==zStateColumn) ? 719:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 34 & r_state==zStateColumn) ? 646:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 36 & r_state==zStateColumn) ? 593:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 38 & r_state==zStateColumn) ? 602:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 40 & r_state==zStateColumn) ? 666:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 42 & r_state==zStateColumn) ? 501:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 44 & r_state==zStateColumn) ? 737:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 46 & r_state==zStateColumn) ? 490:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 48 & r_state==zStateColumn) ? 558:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 50 & r_state==zStateColumn) ? 706:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 52 & r_state==zStateColumn) ? 474:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 54 & r_state==zStateColumn) ? 635:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 56 & r_state==zStateColumn) ? 469:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 58 & r_state==zStateColumn) ? 494:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 60 & r_state==zStateColumn) ? 714:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 62 & r_state==zStateColumn) ? 605:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 64 & r_state==zStateColumn) ? 707:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 66 & r_state==zStateColumn) ? 643:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 68 & r_state==zStateColumn) ? 579:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 70 & r_state==zStateColumn) ? 770:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 72 & r_state==zStateColumn) ? 405:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 74 & r_state==zStateColumn) ? 779:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 76 & r_state==zStateColumn) ? 514:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 78 & r_state==zStateColumn) ? 581:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 80 & r_state==zStateColumn) ? 746:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 82 & r_state==zStateColumn) ? 611:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 84 & r_state==zStateColumn) ? 510:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 86 & r_state==zStateColumn) ? 467:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 88 & r_state==zStateColumn) ? 502:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 90 & r_state==zStateColumn) ? 742:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 92 & r_state==zStateColumn) ? 538:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 94 & r_state==zStateColumn) ? 786:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 96 & r_state==zStateColumn) ? 792:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 98 & r_state==zStateColumn) ? 511:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 100 & r_state==zStateColumn) ? 597:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 102 & r_state==zStateColumn) ? 451:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 104 & r_state==zStateColumn) ? 518:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 106 & r_state==zStateColumn) ? 486:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 108 & r_state==zStateColumn) ? 734:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 110 & r_state==zStateColumn) ? 460:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 112 & r_state==zStateColumn) ? 690:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 114 & r_state==zStateColumn) ? 799:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 116 & r_state==zStateColumn) ? 439:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 118 & r_state==zStateColumn) ? 425:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 120 & r_state==zStateColumn) ? 727:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 122 & r_state==zStateColumn) ? 638:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 124 & r_state==zStateColumn) ? 541:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 126 & r_state==zStateColumn) ? 658:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 128 & r_state==zStateColumn) ? 448:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 130 & r_state==zStateColumn) ? 675:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 132 & r_state==zStateColumn) ? 774:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 134 & r_state==zStateColumn) ? 747:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 136 & r_state==zStateColumn) ? 594:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 138 & r_state==zStateColumn) ? 503:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 140 & r_state==zStateColumn) ? 694:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 142 & r_state==zStateColumn) ? 663:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 144 & r_state==zStateColumn) ? 656:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 146 & r_state==zStateColumn) ? 542:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 148 & r_state==zStateColumn) ? 426:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 150 & r_state==zStateColumn) ? 495:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 152 & r_state==zStateColumn) ? 562:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 154 & r_state==zStateColumn) ? 534:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 156 & r_state==zStateColumn) ? 619:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 158 & r_state==zStateColumn) ? 598:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 160 & r_state==zStateColumn) ? 441:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 162 & r_state==zStateColumn) ? 606:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 164 & r_state==zStateColumn) ? 669:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 166 & r_state==zStateColumn) ? 479:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 168 & r_state==zStateColumn) ? 433:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 170 & r_state==zStateColumn) ? 750:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 172 & r_state==zStateColumn) ? 735:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 174 & r_state==zStateColumn) ? 543:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 176 & r_state==zStateColumn) ? 476:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 178 & r_state==zStateColumn) ? 703:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 180 & r_state==zStateColumn) ? 406:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 182 & r_state==zStateColumn) ? 526:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 184 & r_state==zStateColumn) ? 698:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 186 & r_state==zStateColumn) ? 654:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 188 & r_state==zStateColumn) ? 710:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 190 & r_state==zStateColumn) ? 603:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 192 & r_state==zStateColumn) ? 508:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 194 & r_state==zStateColumn) ? 660:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 196 & r_state==zStateColumn) ? 639:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 198 & r_state==zStateColumn) ? 550:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 200 & r_state==zStateColumn) ? 702:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 202 & r_state==zStateColumn) ? 499:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 204 & r_state==zStateColumn) ? 555:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 206 & r_state==zStateColumn) ? 418:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 208 & r_state==zStateColumn) ? 475:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 210 & r_state==zStateColumn) ? 649:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 212 & r_state==zStateColumn) ? 414:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 214 & r_state==zStateColumn) ? 522:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 216 & r_state==zStateColumn) ? 429:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 218 & r_state==zStateColumn) ? 430:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 220 & r_state==zStateColumn) ? 626:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 222 & r_state==zStateColumn) ? 679:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 224 & r_state==zStateColumn) ? 560:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 226 & r_state==zStateColumn) ? 488:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 228 & r_state==zStateColumn) ? 647:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 230 & r_state==zStateColumn) ? 789:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 232 & r_state==zStateColumn) ? 740:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 234 & r_state==zStateColumn) ? 644:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 236 & r_state==zStateColumn) ? 715:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 238 & r_state==zStateColumn) ? 755:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 240 & r_state==zStateColumn) ? 716:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 242 & r_state==zStateColumn) ? 712:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 244 & r_state==zStateColumn) ? 556:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 246 & r_state==zStateColumn) ? 771:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 248 & r_state==zStateColumn) ? 577:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 250 & r_state==zStateColumn) ? 757:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 252 & r_state==zStateColumn) ? 767:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 254 & r_state==zStateColumn) ? 574:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 256 & r_state==zStateColumn) ? 417:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 258 & r_state==zStateColumn) ? 797:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 260 & r_state==zStateColumn) ? 756:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 262 & r_state==zStateColumn) ? 795:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 264 & r_state==zStateColumn) ? 468:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 266 & r_state==zStateColumn) ? 437:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 268 & r_state==zStateColumn) ? 713:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 270 & r_state==zStateColumn) ? 442:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 272 & r_state==zStateColumn) ? 485:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 274 & r_state==zStateColumn) ? 662:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 276 & r_state==zStateColumn) ? 733:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 278 & r_state==zStateColumn) ? 738:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 280 & r_state==zStateColumn) ? 772:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 282 & r_state==zStateColumn) ? 424:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 284 & r_state==zStateColumn) ? 627:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 286 & r_state==zStateColumn) ? 483:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 288 & r_state==zStateColumn) ? 496:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 290 & r_state==zStateColumn) ? 739:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 292 & r_state==zStateColumn) ? 447:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 294 & r_state==zStateColumn) ? 730:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 296 & r_state==zStateColumn) ? 773:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 298 & r_state==zStateColumn) ? 552:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 300 & r_state==zStateColumn) ? 567:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 302 & r_state==zStateColumn) ? 570:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 304 & r_state==zStateColumn) ? 465:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 306 & r_state==zStateColumn) ? 436:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 308 & r_state==zStateColumn) ? 699:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 310 & r_state==zStateColumn) ? 686:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 312 & r_state==zStateColumn) ? 516:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 314 & r_state==zStateColumn) ? 599:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 316 & r_state==zStateColumn) ? 458:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 318 & r_state==zStateColumn) ? 403:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 320 & r_state==zStateColumn) ? 614:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 322 & r_state==zStateColumn) ? 507:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 324 & r_state==zStateColumn) ? 587:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 326 & r_state==zStateColumn) ? 415:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 328 & r_state==zStateColumn) ? 765:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 330 & r_state==zStateColumn) ? 749:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 332 & r_state==zStateColumn) ? 708:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 334 & r_state==zStateColumn) ? 551:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 336 & r_state==zStateColumn) ? 532:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 338 & r_state==zStateColumn) ? 717:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 340 & r_state==zStateColumn) ? 736:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 342 & r_state==zStateColumn) ? 470:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 344 & r_state==zStateColumn) ? 701:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 346 & r_state==zStateColumn) ? 423:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 348 & r_state==zStateColumn) ? 722:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 350 & r_state==zStateColumn) ? 410:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 352 & r_state==zStateColumn) ? 412:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 354 & r_state==zStateColumn) ? 684:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 356 & r_state==zStateColumn) ? 407:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 358 & r_state==zStateColumn) ? 762:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 360 & r_state==zStateColumn) ? 493:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 362 & r_state==zStateColumn) ? 631:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 364 & r_state==zStateColumn) ? 731:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 366 & r_state==zStateColumn) ? 623:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 368 & r_state==zStateColumn) ? 629:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 370 & r_state==zStateColumn) ? 709:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 372 & r_state==zStateColumn) ? 536:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 374 & r_state==zStateColumn) ? 787:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 376 & r_state==zStateColumn) ? 440:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 378 & r_state==zStateColumn) ? 677:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 380 & r_state==zStateColumn) ? 705:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 382 & r_state==zStateColumn) ? 650:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 384 & r_state==zStateColumn) ? 726:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 386 & r_state==zStateColumn) ? 798:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 388 & r_state==zStateColumn) ? 785:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 390 & r_state==zStateColumn) ? 758:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 392 & r_state==zStateColumn) ? 784:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 394 & r_state==zStateColumn) ? 793:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 396 & r_state==zStateColumn) ? 601:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 398 & r_state==zStateColumn) ? 461:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 400 & r_state==zStateColumn) ? 732:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 402 & r_state==zStateColumn) ? 512:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 404 & r_state==zStateColumn) ? 636:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 406 & r_state==zStateColumn) ? 563:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 408 & r_state==zStateColumn) ? 664:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 410 & r_state==zStateColumn) ? 620:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 412 & r_state==zStateColumn) ? 416:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 414 & r_state==zStateColumn) ? 763:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 416 & r_state==zStateColumn) ? 464:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 418 & r_state==zStateColumn) ? 420:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 420 & r_state==zStateColumn) ? 788:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 422 & r_state==zStateColumn) ? 427:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 424 & r_state==zStateColumn) ? 604:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 426 & r_state==zStateColumn) ? 624:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 428 & r_state==zStateColumn) ? 431:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 430 & r_state==zStateColumn) ? 681:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 432 & r_state==zStateColumn) ? 472:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 434 & r_state==zStateColumn) ? 572:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 436 & r_state==zStateColumn) ? 776:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 438 & r_state==zStateColumn) ? 751:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 440 & r_state==zStateColumn) ? 408:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 442 & r_state==zStateColumn) ? 676:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 444 & r_state==zStateColumn) ? 582:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 446 & r_state==zStateColumn) ? 782:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 448 & r_state==zStateColumn) ? 724:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 450 & r_state==zStateColumn) ? 688:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 452 & r_state==zStateColumn) ? 704:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 454 & r_state==zStateColumn) ? 595:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 456 & r_state==zStateColumn) ? 689:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 458 & r_state==zStateColumn) ? 584:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 460 & r_state==zStateColumn) ? 487:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 462 & r_state==zStateColumn) ? 531:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 464 & r_state==zStateColumn) ? 564:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 466 & r_state==zStateColumn) ? 553:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 468 & r_state==zStateColumn) ? 540:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 470 & r_state==zStateColumn) ? 759:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 472 & r_state==zStateColumn) ? 504:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 474 & r_state==zStateColumn) ? 668:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 476 & r_state==zStateColumn) ? 497:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 478 & r_state==zStateColumn) ? 443:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 480 & r_state==zStateColumn) ? 696:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 482 & r_state==zStateColumn) ? 600:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 484 & r_state==zStateColumn) ? 764:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 486 & r_state==zStateColumn) ? 723:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 488 & r_state==zStateColumn) ? 428:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 490 & r_state==zStateColumn) ? 725:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 492 & r_state==zStateColumn) ? 576:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 494 & r_state==zStateColumn) ? 670:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 496 & r_state==zStateColumn) ? 492:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 498 & r_state==zStateColumn) ? 632:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 500 & r_state==zStateColumn) ? 432:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 502 & r_state==zStateColumn) ? 462:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 504 & r_state==zStateColumn) ? 672:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 506 & r_state==zStateColumn) ? 768:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 508 & r_state==zStateColumn) ? 590:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 510 & r_state==zStateColumn) ? 790:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 512 & r_state==zStateColumn) ? 752:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 514 & r_state==zStateColumn) ? 528:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 516 & r_state==zStateColumn) ? 728:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 518 & r_state==zStateColumn) ? 667:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 520 & r_state==zStateColumn) ? 608:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 522 & r_state==zStateColumn) ? 748:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 524 & r_state==zStateColumn) ? 456:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 526 & r_state==zStateColumn) ? 655:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 528 & r_state==zStateColumn) ? 753:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 530 & r_state==zStateColumn) ? 529:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 532 & r_state==zStateColumn) ? 665:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 534 & r_state==zStateColumn) ? 583:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 536 & r_state==zStateColumn) ? 625:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 538 & r_state==zStateColumn) ? 700:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 540 & r_state==zStateColumn) ? 513:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 542 & r_state==zStateColumn) ? 471:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 544 & r_state==zStateColumn) ? 400:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 546 & r_state==zStateColumn) ? 769:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 548 & r_state==zStateColumn) ? 548:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 550 & r_state==zStateColumn) ? 691:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 552 & r_state==zStateColumn) ? 524:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 554 & r_state==zStateColumn) ? 473:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 556 & r_state==zStateColumn) ? 612:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 558 & r_state==zStateColumn) ? 671:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 560 & r_state==zStateColumn) ? 409:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 562 & r_state==zStateColumn) ? 796:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 564 & r_state==zStateColumn) ? 640:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 566 & r_state==zStateColumn) ? 459:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 568 & r_state==zStateColumn) ? 498:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 570 & r_state==zStateColumn) ? 744:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 572 & r_state==zStateColumn) ? 449:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 574 & r_state==zStateColumn) ? 783:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 576 & r_state==zStateColumn) ? 777:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 578 & r_state==zStateColumn) ? 621:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 580 & r_state==zStateColumn) ? 743:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 582 & r_state==zStateColumn) ? 547:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 584 & r_state==zStateColumn) ? 680:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 586 & r_state==zStateColumn) ? 505:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 588 & r_state==zStateColumn) ? 480:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 590 & r_state==zStateColumn) ? 463:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 592 & r_state==zStateColumn) ? 444:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 594 & r_state==zStateColumn) ? 500:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 596 & r_state==zStateColumn) ? 745:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 598 & r_state==zStateColumn) ? 575:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 600 & r_state==zStateColumn) ? 457:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 602 & r_state==zStateColumn) ? 729:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 604 & r_state==zStateColumn) ? 673:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 606 & r_state==zStateColumn) ? 711:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 608 & r_state==zStateColumn) ? 648:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 610 & r_state==zStateColumn) ? 549:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 612 & r_state==zStateColumn) ? 533:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 614 & r_state==zStateColumn) ? 535:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 616 & r_state==zStateColumn) ? 780:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 618 & r_state==zStateColumn) ? 445:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 620 & r_state==zStateColumn) ? 435:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 622 & r_state==zStateColumn) ? 454:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 624 & r_state==zStateColumn) ? 718:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 626 & r_state==zStateColumn) ? 674:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 628 & r_state==zStateColumn) ? 580:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 630 & r_state==zStateColumn) ? 659:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 632 & r_state==zStateColumn) ? 544:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 634 & r_state==zStateColumn) ? 484:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 636 & r_state==zStateColumn) ? 628:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 638 & r_state==zStateColumn) ? 519:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 640 & r_state==zStateColumn) ? 609:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 642 & r_state==zStateColumn) ? 645:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 644 & r_state==zStateColumn) ? 692:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 646 & r_state==zStateColumn) ? 791:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 648 & r_state==zStateColumn) ? 413:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 650 & r_state==zStateColumn) ? 585:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 652 & r_state==zStateColumn) ? 661:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 654 & r_state==zStateColumn) ? 687:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 656 & r_state==zStateColumn) ? 450:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 658 & r_state==zStateColumn) ? 452:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 660 & r_state==zStateColumn) ? 633:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 662 & r_state==zStateColumn) ? 559:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 664 & r_state==zStateColumn) ? 720:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 666 & r_state==zStateColumn) ? 401:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 668 & r_state==zStateColumn) ? 481:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 670 & r_state==zStateColumn) ? 515:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 672 & r_state==zStateColumn) ? 634:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 674 & r_state==zStateColumn) ? 721:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 676 & r_state==zStateColumn) ? 568:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 678 & r_state==zStateColumn) ? 527:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 680 & r_state==zStateColumn) ? 588:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 682 & r_state==zStateColumn) ? 610:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 684 & r_state==zStateColumn) ? 545:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 686 & r_state==zStateColumn) ? 419:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 688 & r_state==zStateColumn) ? 569:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 690 & r_state==zStateColumn) ? 778:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 692 & r_state==zStateColumn) ? 754:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 694 & r_state==zStateColumn) ? 775:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 696 & r_state==zStateColumn) ? 477:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 698 & r_state==zStateColumn) ? 546:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 700 & r_state==zStateColumn) ? 586:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 702 & r_state==zStateColumn) ? 607:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 704 & r_state==zStateColumn) ? 613:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 706 & r_state==zStateColumn) ? 652:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 708 & r_state==zStateColumn) ? 622:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 710 & r_state==zStateColumn) ? 571:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 712 & r_state==zStateColumn) ? 592:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 714 & r_state==zStateColumn) ? 760:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 716 & r_state==zStateColumn) ? 630:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 718 & r_state==zStateColumn) ? 491:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 720 & r_state==zStateColumn) ? 557:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 722 & r_state==zStateColumn) ? 693:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 724 & r_state==zStateColumn) ? 637:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 726 & r_state==zStateColumn) ? 695:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 728 & r_state==zStateColumn) ? 596:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 730 & r_state==zStateColumn) ? 616:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 732 & r_state==zStateColumn) ? 520:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 734 & r_state==zStateColumn) ? 411:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 736 & r_state==zStateColumn) ? 578:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 738 & r_state==zStateColumn) ? 617:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 740 & r_state==zStateColumn) ? 641:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 742 & r_state==zStateColumn) ? 523:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 744 & r_state==zStateColumn) ? 446:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 746 & r_state==zStateColumn) ? 685:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 748 & r_state==zStateColumn) ? 741:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 750 & r_state==zStateColumn) ? 682:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 752 & r_state==zStateColumn) ? 402:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 754 & r_state==zStateColumn) ? 697:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 756 & r_state==zStateColumn) ? 466:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 758 & r_state==zStateColumn) ? 615:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 760 & r_state==zStateColumn) ? 521:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 762 & r_state==zStateColumn) ? 573:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 764 & r_state==zStateColumn) ? 506:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 766 & r_state==zStateColumn) ? 683:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 768 & r_state==zStateColumn) ? 781:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 770 & r_state==zStateColumn) ? 530:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 772 & r_state==zStateColumn) ? 589:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 774 & r_state==zStateColumn) ? 591:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 776 & r_state==zStateColumn) ? 525:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 778 & r_state==zStateColumn) ? 761:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 780 & r_state==zStateColumn) ? 618:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 782 & r_state==zStateColumn) ? 651:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 784 & r_state==zStateColumn) ? 478:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 786 & r_state==zStateColumn) ? 482:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 788 & r_state==zStateColumn) ? 438:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 790 & r_state==zStateColumn) ? 539:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 792 & r_state==zStateColumn) ? 421:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 794 & r_state==zStateColumn) ? 453:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 796 & r_state==zStateColumn) ? 653:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 798 & r_state==zStateColumn) ? 455:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 800 & r_state==zStateColumn) ? 272:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 802 & r_state==zStateColumn) ? 333:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 804 & r_state==zStateColumn) ? 376:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 806 & r_state==zStateColumn) ? 159:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 808 & r_state==zStateColumn) ? 5:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 810 & r_state==zStateColumn) ? 36:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 812 & r_state==zStateColumn) ? 90:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 814 & r_state==zStateColumn) ? 178:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 816 & r_state==zStateColumn) ? 220:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 818 & r_state==zStateColumn) ? 280:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 820 & r_state==zStateColumn) ? 175:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 822 & r_state==zStateColumn) ? 367:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 824 & r_state==zStateColumn) ? 176:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 826 & r_state==zStateColumn) ? 324:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 828 & r_state==zStateColumn) ? 106:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 830 & r_state==zStateColumn) ? 163:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 832 & r_state==zStateColumn) ? 206:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 834 & r_state==zStateColumn) ? 128:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 836 & r_state==zStateColumn) ? 103:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 838 & r_state==zStateColumn) ? 343:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 840 & r_state==zStateColumn) ? 209:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 842 & r_state==zStateColumn) ? 396:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 844 & r_state==zStateColumn) ? 7:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 846 & r_state==zStateColumn) ? 173:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 848 & r_state==zStateColumn) ? 141:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 850 & r_state==zStateColumn) ? 59:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 852 & r_state==zStateColumn) ? 74:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 854 & r_state==zStateColumn) ? 211:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 856 & r_state==zStateColumn) ? 244:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 858 & r_state==zStateColumn) ? 108:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 860 & r_state==zStateColumn) ? 109:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 862 & r_state==zStateColumn) ? 214:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 864 & r_state==zStateColumn) ? 250:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 866 & r_state==zStateColumn) ? 84:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 868 & r_state==zStateColumn) ? 10:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 870 & r_state==zStateColumn) ? 310:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 872 & r_state==zStateColumn) ? 153:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 874 & r_state==zStateColumn) ? 133:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 876 & r_state==zStateColumn) ? 394:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 878 & r_state==zStateColumn) ? 58:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 880 & r_state==zStateColumn) ? 188:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 882 & r_state==zStateColumn) ? 80:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 884 & r_state==zStateColumn) ? 135:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 886 & r_state==zStateColumn) ? 239:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 888 & r_state==zStateColumn) ? 296:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 890 & r_state==zStateColumn) ? 309:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 892 & r_state==zStateColumn) ? 372:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 894 & r_state==zStateColumn) ? 146:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 896 & r_state==zStateColumn) ? 64:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 898 & r_state==zStateColumn) ? 286:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 900 & r_state==zStateColumn) ? 328:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 902 & r_state==zStateColumn) ? 51:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 904 & r_state==zStateColumn) ? 329:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 906 & r_state==zStateColumn) ? 397:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 908 & r_state==zStateColumn) ? 311:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 910 & r_state==zStateColumn) ? 399:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 912 & r_state==zStateColumn) ? 262:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 914 & r_state==zStateColumn) ? 300:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 916 & r_state==zStateColumn) ? 158:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 918 & r_state==zStateColumn) ? 283:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 920 & r_state==zStateColumn) ? 55:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 922 & r_state==zStateColumn) ? 199:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 924 & r_state==zStateColumn) ? 251:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 926 & r_state==zStateColumn) ? 295:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 928 & r_state==zStateColumn) ? 208:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 930 & r_state==zStateColumn) ? 152:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 932 & r_state==zStateColumn) ? 378:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 934 & r_state==zStateColumn) ? 43:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 936 & r_state==zStateColumn) ? 132:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 938 & r_state==zStateColumn) ? 28:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 940 & r_state==zStateColumn) ? 171:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 942 & r_state==zStateColumn) ? 271:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 944 & r_state==zStateColumn) ? 216:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 946 & r_state==zStateColumn) ? 277:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 948 & r_state==zStateColumn) ? 26:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 950 & r_state==zStateColumn) ? 104:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 952 & r_state==zStateColumn) ? 88:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 954 & r_state==zStateColumn) ? 348:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 956 & r_state==zStateColumn) ? 392:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 958 & r_state==zStateColumn) ? 83:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 960 & r_state==zStateColumn) ? 294:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 962 & r_state==zStateColumn) ? 334:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 964 & r_state==zStateColumn) ? 393:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 966 & r_state==zStateColumn) ? 143:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 968 & r_state==zStateColumn) ? 317:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 970 & r_state==zStateColumn) ? 136:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 972 & r_state==zStateColumn) ? 53:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 974 & r_state==zStateColumn) ? 230:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 976 & r_state==zStateColumn) ? 113:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 978 & r_state==zStateColumn) ? 2:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 980 & r_state==zStateColumn) ? 23:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 982 & r_state==zStateColumn) ? 359:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 984 & r_state==zStateColumn) ? 248:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 986 & r_state==zStateColumn) ? 180:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 988 & r_state==zStateColumn) ? 29:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 990 & r_state==zStateColumn) ? 75:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 992 & r_state==zStateColumn) ? 144:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 994 & r_state==zStateColumn) ? 238:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 996 & r_state==zStateColumn) ? 284:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 998 & r_state==zStateColumn) ? 101:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1000 & r_state==zStateColumn) ? 297:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1002 & r_state==zStateColumn) ? 21:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1004 & r_state==zStateColumn) ? 44:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1006 & r_state==zStateColumn) ? 69:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1008 & r_state==zStateColumn) ? 236:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1010 & r_state==zStateColumn) ? 293:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1012 & r_state==zStateColumn) ? 382:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1014 & r_state==zStateColumn) ? 161:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1016 & r_state==zStateColumn) ? 96:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1018 & r_state==zStateColumn) ? 6:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1020 & r_state==zStateColumn) ? 42:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1022 & r_state==zStateColumn) ? 49:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1024 & r_state==zStateColumn) ? 201:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1026 & r_state==zStateColumn) ? 270:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1028 & r_state==zStateColumn) ? 38:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1030 & r_state==zStateColumn) ? 335:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1032 & r_state==zStateColumn) ? 156:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1034 & r_state==zStateColumn) ? 12:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1036 & r_state==zStateColumn) ? 52:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1038 & r_state==zStateColumn) ? 319:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1040 & r_state==zStateColumn) ? 366:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1042 & r_state==zStateColumn) ? 380:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1044 & r_state==zStateColumn) ? 107:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1046 & r_state==zStateColumn) ? 371:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1048 & r_state==zStateColumn) ? 276:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1050 & r_state==zStateColumn) ? 388:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1052 & r_state==zStateColumn) ? 91:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1054 & r_state==zStateColumn) ? 339:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1056 & r_state==zStateColumn) ? 257:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1058 & r_state==zStateColumn) ? 265:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1060 & r_state==zStateColumn) ? 385:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1062 & r_state==zStateColumn) ? 231:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1064 & r_state==zStateColumn) ? 168:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1066 & r_state==zStateColumn) ? 306:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1068 & r_state==zStateColumn) ? 77:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1070 & r_state==zStateColumn) ? 307:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1072 & r_state==zStateColumn) ? 186:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1074 & r_state==zStateColumn) ? 13:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1076 & r_state==zStateColumn) ? 46:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1078 & r_state==zStateColumn) ? 395:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1080 & r_state==zStateColumn) ? 234:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1082 & r_state==zStateColumn) ? 62:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1084 & r_state==zStateColumn) ? 73:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1086 & r_state==zStateColumn) ? 87:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1088 & r_state==zStateColumn) ? 316:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1090 & r_state==zStateColumn) ? 342:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1092 & r_state==zStateColumn) ? 349:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1094 & r_state==zStateColumn) ? 291:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1096 & r_state==zStateColumn) ? 274:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1098 & r_state==zStateColumn) ? 305:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1100 & r_state==zStateColumn) ? 99:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1102 & r_state==zStateColumn) ? 167:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1104 & r_state==zStateColumn) ? 149:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1106 & r_state==zStateColumn) ? 233:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1108 & r_state==zStateColumn) ? 14:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1110 & r_state==zStateColumn) ? 102:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1112 & r_state==zStateColumn) ? 122:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1114 & r_state==zStateColumn) ? 360:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1116 & r_state==zStateColumn) ? 24:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1118 & r_state==zStateColumn) ? 331:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1120 & r_state==zStateColumn) ? 112:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1122 & r_state==zStateColumn) ? 9:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1124 & r_state==zStateColumn) ? 76:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1126 & r_state==zStateColumn) ? 203:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1128 & r_state==zStateColumn) ? 232:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1130 & r_state==zStateColumn) ? 0:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1132 & r_state==zStateColumn) ? 1:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1134 & r_state==zStateColumn) ? 150:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1136 & r_state==zStateColumn) ? 338:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1138 & r_state==zStateColumn) ? 344:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1140 & r_state==zStateColumn) ? 151:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1142 & r_state==zStateColumn) ? 355:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1144 & r_state==zStateColumn) ? 217:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1146 & r_state==zStateColumn) ? 381:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1148 & r_state==zStateColumn) ? 127:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1150 & r_state==zStateColumn) ? 299:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1152 & r_state==zStateColumn) ? 246:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1154 & r_state==zStateColumn) ? 124:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1156 & r_state==zStateColumn) ? 368:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1158 & r_state==zStateColumn) ? 34:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1160 & r_state==zStateColumn) ? 314:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1162 & r_state==zStateColumn) ? 39:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1164 & r_state==zStateColumn) ? 222:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1166 & r_state==zStateColumn) ? 267:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1168 & r_state==zStateColumn) ? 229:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1170 & r_state==zStateColumn) ? 325:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1172 & r_state==zStateColumn) ? 350:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1174 & r_state==zStateColumn) ? 162:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1176 & r_state==zStateColumn) ? 340:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1178 & r_state==zStateColumn) ? 386:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1180 & r_state==zStateColumn) ? 254:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1182 & r_state==zStateColumn) ? 387:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1184 & r_state==zStateColumn) ? 356:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1186 & r_state==zStateColumn) ? 18:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1188 & r_state==zStateColumn) ? 68:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1190 & r_state==zStateColumn) ? 227:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1192 & r_state==zStateColumn) ? 364:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1194 & r_state==zStateColumn) ? 50:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1196 & r_state==zStateColumn) ? 79:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1198 & r_state==zStateColumn) ? 157:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1200 & r_state==zStateColumn) ? 241:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1202 & r_state==zStateColumn) ? 198:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1204 & r_state==zStateColumn) ? 19:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1206 & r_state==zStateColumn) ? 95:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1208 & r_state==zStateColumn) ? 212:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1210 & r_state==zStateColumn) ? 31:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1212 & r_state==zStateColumn) ? 81:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1214 & r_state==zStateColumn) ? 351:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1216 & r_state==zStateColumn) ? 260:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1218 & r_state==zStateColumn) ? 320:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1220 & r_state==zStateColumn) ? 341:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1222 & r_state==zStateColumn) ? 41:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1224 & r_state==zStateColumn) ? 278:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1226 & r_state==zStateColumn) ? 352:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1228 & r_state==zStateColumn) ? 160:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1230 & r_state==zStateColumn) ? 379:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1232 & r_state==zStateColumn) ? 365:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1234 & r_state==zStateColumn) ? 369:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1236 & r_state==zStateColumn) ? 390:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1238 & r_state==zStateColumn) ? 78:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1240 & r_state==zStateColumn) ? 205:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1242 & r_state==zStateColumn) ? 289:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1244 & r_state==zStateColumn) ? 354:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1246 & r_state==zStateColumn) ? 183:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1248 & r_state==zStateColumn) ? 213:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1250 & r_state==zStateColumn) ? 268:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1252 & r_state==zStateColumn) ? 110:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1254 & r_state==zStateColumn) ? 142:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1256 & r_state==zStateColumn) ? 318:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1258 & r_state==zStateColumn) ? 184:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1260 & r_state==zStateColumn) ? 358:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1262 & r_state==zStateColumn) ? 181:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1264 & r_state==zStateColumn) ? 249:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1266 & r_state==zStateColumn) ? 330:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1268 & r_state==zStateColumn) ? 336:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1270 & r_state==zStateColumn) ? 27:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1272 & r_state==zStateColumn) ? 202:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1274 & r_state==zStateColumn) ? 362:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1276 & r_state==zStateColumn) ? 61:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1278 & r_state==zStateColumn) ? 98:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1280 & r_state==zStateColumn) ? 282:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1282 & r_state==zStateColumn) ? 370:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1284 & r_state==zStateColumn) ? 8:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1286 & r_state==zStateColumn) ? 33:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1288 & r_state==zStateColumn) ? 117:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1290 & r_state==zStateColumn) ? 321:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1292 & r_state==zStateColumn) ? 17:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1294 & r_state==zStateColumn) ? 114:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1296 & r_state==zStateColumn) ? 304:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1298 & r_state==zStateColumn) ? 105:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1300 & r_state==zStateColumn) ? 191:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1302 & r_state==zStateColumn) ? 391:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1304 & r_state==zStateColumn) ? 353:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1306 & r_state==zStateColumn) ? 398:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1308 & r_state==zStateColumn) ? 93:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1310 & r_state==zStateColumn) ? 263:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1312 & r_state==zStateColumn) ? 72:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1314 & r_state==zStateColumn) ? 11:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1316 & r_state==zStateColumn) ? 63:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1318 & r_state==zStateColumn) ? 315:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1320 & r_state==zStateColumn) ? 97:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1322 & r_state==zStateColumn) ? 326:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1324 & r_state==zStateColumn) ? 137:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1326 & r_state==zStateColumn) ? 71:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1328 & r_state==zStateColumn) ? 204:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1330 & r_state==zStateColumn) ? 266:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1332 & r_state==zStateColumn) ? 20:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1334 & r_state==zStateColumn) ? 259:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1336 & r_state==zStateColumn) ? 237:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1338 & r_state==zStateColumn) ? 82:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1340 & r_state==zStateColumn) ? 247:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1342 & r_state==zStateColumn) ? 279:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1344 & r_state==zStateColumn) ? 252:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1346 & r_state==zStateColumn) ? 302:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1348 & r_state==zStateColumn) ? 313:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1350 & r_state==zStateColumn) ? 65:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1352 & r_state==zStateColumn) ? 221:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1354 & r_state==zStateColumn) ? 189:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1356 & r_state==zStateColumn) ? 3:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1358 & r_state==zStateColumn) ? 111:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1360 & r_state==zStateColumn) ? 292:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1362 & r_state==zStateColumn) ? 215:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1364 & r_state==zStateColumn) ? 375:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1366 & r_state==zStateColumn) ? 383:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1368 & r_state==zStateColumn) ? 177:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1370 & r_state==zStateColumn) ? 373:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1372 & r_state==zStateColumn) ? 155:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1374 & r_state==zStateColumn) ? 327:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1376 & r_state==zStateColumn) ? 225:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1378 & r_state==zStateColumn) ? 228:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1380 & r_state==zStateColumn) ? 56:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1382 & r_state==zStateColumn) ? 275:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1384 & r_state==zStateColumn) ? 322:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1386 & r_state==zStateColumn) ? 361:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1388 & r_state==zStateColumn) ? 70:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1390 & r_state==zStateColumn) ? 363:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1392 & r_state==zStateColumn) ? 240:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1394 & r_state==zStateColumn) ? 377:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1396 & r_state==zStateColumn) ? 92:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1398 & r_state==zStateColumn) ? 154:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1400 & r_state==zStateColumn) ? 269:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1402 & r_state==zStateColumn) ? 172:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1404 & r_state==zStateColumn) ? 100:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1406 & r_state==zStateColumn) ? 89:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1408 & r_state==zStateColumn) ? 226:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1410 & r_state==zStateColumn) ? 190:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1412 & r_state==zStateColumn) ? 25:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1414 & r_state==zStateColumn) ? 32:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1416 & r_state==zStateColumn) ? 166:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1418 & r_state==zStateColumn) ? 185:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1420 & r_state==zStateColumn) ? 94:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1422 & r_state==zStateColumn) ? 303:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1424 & r_state==zStateColumn) ? 121:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1426 & r_state==zStateColumn) ? 134:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1428 & r_state==zStateColumn) ? 30:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1430 & r_state==zStateColumn) ? 118:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1432 & r_state==zStateColumn) ? 120:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1434 & r_state==zStateColumn) ? 169:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1436 & r_state==zStateColumn) ? 312:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1438 & r_state==zStateColumn) ? 16:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1440 & r_state==zStateColumn) ? 332:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1442 & r_state==zStateColumn) ? 337:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1444 & r_state==zStateColumn) ? 174:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1446 & r_state==zStateColumn) ? 243:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1448 & r_state==zStateColumn) ? 224:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1450 & r_state==zStateColumn) ? 245:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1452 & r_state==zStateColumn) ? 192:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1454 & r_state==zStateColumn) ? 60:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1456 & r_state==zStateColumn) ? 258:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1458 & r_state==zStateColumn) ? 301:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1460 & r_state==zStateColumn) ? 147:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1462 & r_state==zStateColumn) ? 182:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1464 & r_state==zStateColumn) ? 200:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1466 & r_state==zStateColumn) ? 138:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1468 & r_state==zStateColumn) ? 54:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1470 & r_state==zStateColumn) ? 86:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1472 & r_state==zStateColumn) ? 170:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1474 & r_state==zStateColumn) ? 22:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1476 & r_state==zStateColumn) ? 139:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1478 & r_state==zStateColumn) ? 145:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1480 & r_state==zStateColumn) ? 116:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1482 & r_state==zStateColumn) ? 374:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1484 & r_state==zStateColumn) ? 45:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1486 & r_state==zStateColumn) ? 290:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1488 & r_state==zStateColumn) ? 285:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1490 & r_state==zStateColumn) ? 298:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1492 & r_state==zStateColumn) ? 40:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1494 & r_state==zStateColumn) ? 67:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1496 & r_state==zStateColumn) ? 261:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1498 & r_state==zStateColumn) ? 165:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1500 & r_state==zStateColumn) ? 85:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1502 & r_state==zStateColumn) ? 219:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1504 & r_state==zStateColumn) ? 256:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1506 & r_state==zStateColumn) ? 264:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1508 & r_state==zStateColumn) ? 346:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1510 & r_state==zStateColumn) ? 119:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1512 & r_state==zStateColumn) ? 130:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1514 & r_state==zStateColumn) ? 125:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1516 & r_state==zStateColumn) ? 195:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1518 & r_state==zStateColumn) ? 235:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1520 & r_state==zStateColumn) ? 357:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1522 & r_state==zStateColumn) ? 389:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1524 & r_state==zStateColumn) ? 179:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1526 & r_state==zStateColumn) ? 207:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1528 & r_state==zStateColumn) ? 242:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1530 & r_state==zStateColumn) ? 164:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1532 & r_state==zStateColumn) ? 15:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1534 & r_state==zStateColumn) ? 126:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1536 & r_state==zStateColumn) ? 253:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1538 & r_state==zStateColumn) ? 273:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1540 & r_state==zStateColumn) ? 35:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1542 & r_state==zStateColumn) ? 123:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1544 & r_state==zStateColumn) ? 140:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1546 & r_state==zStateColumn) ? 148:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1548 & r_state==zStateColumn) ? 66:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1550 & r_state==zStateColumn) ? 347:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1552 & r_state==zStateColumn) ? 218:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1554 & r_state==zStateColumn) ? 288:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1556 & r_state==zStateColumn) ? 345:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1558 & r_state==zStateColumn) ? 37:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1560 & r_state==zStateColumn) ? 308:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1562 & r_state==zStateColumn) ? 384:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1564 & r_state==zStateColumn) ? 223:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1566 & r_state==zStateColumn) ? 287:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1568 & r_state==zStateColumn) ? 196:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1570 & r_state==zStateColumn) ? 194:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1572 & r_state==zStateColumn) ? 47:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1574 & r_state==zStateColumn) ? 187:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1576 & r_state==zStateColumn) ? 210:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1578 & r_state==zStateColumn) ? 115:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1580 & r_state==zStateColumn) ? 255:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1582 & r_state==zStateColumn) ? 323:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1584 & r_state==zStateColumn) ? 48:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1586 & r_state==zStateColumn) ? 197:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1588 & r_state==zStateColumn) ? 4:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1590 & r_state==zStateColumn) ? 131:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1592 & r_state==zStateColumn) ? 281:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1594 & r_state==zStateColumn) ? 129:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1596 & r_state==zStateColumn) ? 193:
			/**/
			/**/
		        /**/
			/**/
		        /**/ 
			(r_counter == 1598 & r_state==zStateColumn) ? 57:
			/**/
			/**/
		        /**/
			/**/
			/**/
			 /**/
			(r_counter == 0 & r_state==zStateEstimate) ? 196:
			/**/
			/**/
			 /**/
			(r_counter == 1 & r_state==zStateEstimate) ? 784:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 3 & r_state==zStateEstimate) ? 140:
			/**/
			/**/
			 /**/
			(r_counter == 4 & r_state==zStateEstimate) ? 772:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 6 & r_state==zStateEstimate) ? 200:
			/**/
			/**/
			 /**/
			(r_counter == 7 & r_state==zStateEstimate) ? 732:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 9 & r_state==zStateEstimate) ? 201:
			/**/
			/**/
			 /**/
			(r_counter == 10 & r_state==zStateEstimate) ? 512:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 12 & r_state==zStateEstimate) ? 202:
			/**/
			/**/
			 /**/
			(r_counter == 13 & r_state==zStateEstimate) ? 636:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 15 & r_state==zStateEstimate) ? 112:
			/**/
			/**/
			 /**/
			(r_counter == 16 & r_state==zStateEstimate) ? 560:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 18 & r_state==zStateEstimate) ? 204:
			/**/
			/**/
			 /**/
			(r_counter == 19 & r_state==zStateEstimate) ? 664:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 21 & r_state==zStateEstimate) ? 205:
			/**/
			/**/
			 /**/
			(r_counter == 22 & r_state==zStateEstimate) ? 620:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 24 & r_state==zStateEstimate) ? 206:
			/**/
			/**/
			 /**/
			(r_counter == 25 & r_state==zStateEstimate) ? 416:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 27 & r_state==zStateEstimate) ? 48:
			/**/
			/**/
			 /**/
			(r_counter == 28 & r_state==zStateEstimate) ? 792:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 30 & r_state==zStateEstimate) ? 208:
			/**/
			/**/
			 /**/
			(r_counter == 31 & r_state==zStateEstimate) ? 464:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 33 & r_state==zStateEstimate) ? 209:
			/**/
			/**/
			 /**/
			(r_counter == 34 & r_state==zStateEstimate) ? 420:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 36 & r_state==zStateEstimate) ? 210:
			/**/
			/**/
			 /**/
			(r_counter == 37 & r_state==zStateEstimate) ? 788:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 39 & r_state==zStateEstimate) ? 88:
			/**/
			/**/
			 /**/
			(r_counter == 40 & r_state==zStateEstimate) ? 476:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 42 & r_state==zStateEstimate) ? 212:
			/**/
			/**/
			 /**/
			(r_counter == 43 & r_state==zStateEstimate) ? 604:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 45 & r_state==zStateEstimate) ? 213:
			/**/
			/**/
			 /**/
			(r_counter == 46 & r_state==zStateEstimate) ? 624:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 48 & r_state==zStateEstimate) ? 144:
			/**/
			/**/
			 /**/
			(r_counter == 49 & r_state==zStateEstimate) ? 496:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 51 & r_state==zStateEstimate) ? 116:
			/**/
			/**/
			 /**/
			(r_counter == 52 & r_state==zStateEstimate) ? 740:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 54 & r_state==zStateEstimate) ? 216:
			/**/
			/**/
			 /**/
			(r_counter == 55 & r_state==zStateEstimate) ? 472:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 57 & r_state==zStateEstimate) ? 217:
			/**/
			/**/
			 /**/
			(r_counter == 58 & r_state==zStateEstimate) ? 572:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 60 & r_state==zStateEstimate) ? 218:
			/**/
			/**/
			 /**/
			(r_counter == 61 & r_state==zStateEstimate) ? 776:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 63 & r_state==zStateEstimate) ? 117:
			/**/
			/**/
			 /**/
			(r_counter == 64 & r_state==zStateEstimate) ? 644:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 66 & r_state==zStateEstimate) ? 220:
			/**/
			/**/
			 /**/
			(r_counter == 67 & r_state==zStateEstimate) ? 408:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 69 & r_state==zStateEstimate) ? 148:
			/**/
			/**/
			 /**/
			(r_counter == 70 & r_state==zStateEstimate) ? 773:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 72 & r_state==zStateEstimate) ? 221:
			/**/
			/**/
			 /**/
			(r_counter == 73 & r_state==zStateEstimate) ? 676:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 75 & r_state==zStateEstimate) ? 149:
			/**/
			/**/
			 /**/
			(r_counter == 76 & r_state==zStateEstimate) ? 552:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 78 & r_state==zStateEstimate) ? 224:
			/**/
			/**/
			 /**/
			(r_counter == 79 & r_state==zStateEstimate) ? 724:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 81 & r_state==zStateEstimate) ? 225:
			/**/
			/**/
			 /**/
			(r_counter == 82 & r_state==zStateEstimate) ? 688:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 84 & r_state==zStateEstimate) ? 226:
			/**/
			/**/
			 /**/
			(r_counter == 85 & r_state==zStateEstimate) ? 704:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 87 & r_state==zStateEstimate) ? 72:
			/**/
			/**/
			 /**/
			(r_counter == 88 & r_state==zStateEstimate) ? 656:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 90 & r_state==zStateEstimate) ? 152:
			/**/
			/**/
			 /**/
			(r_counter == 91 & r_state==zStateEstimate) ? 465:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 93 & r_state==zStateEstimate) ? 228:
			/**/
			/**/
			 /**/
			(r_counter == 94 & r_state==zStateEstimate) ? 689:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 96 & r_state==zStateEstimate) ? 229:
			/**/
			/**/
			 /**/
			(r_counter == 97 & r_state==zStateEstimate) ? 584:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 99 & r_state==zStateEstimate) ? 120:
			/**/
			/**/
			 /**/
			(r_counter == 100 & r_state==zStateEstimate) ? 716:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 102 & r_state==zStateEstimate) ? 232:
			/**/
			/**/
			 /**/
			(r_counter == 103 & r_state==zStateEstimate) ? 564:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 105 & r_state==zStateEstimate) ? 233:
			/**/
			/**/
			 /**/
			(r_counter == 106 & r_state==zStateEstimate) ? 553:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 108 & r_state==zStateEstimate) ? 234:
			/**/
			/**/
			 /**/
			(r_counter == 109 & r_state==zStateEstimate) ? 540:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 111 & r_state==zStateEstimate) ? 153:
			/**/
			/**/
			 /**/
			(r_counter == 112 & r_state==zStateEstimate) ? 436:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 114 & r_state==zStateEstimate) ? 236:
			/**/
			/**/
			 /**/
			(r_counter == 115 & r_state==zStateEstimate) ? 504:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 117 & r_state==zStateEstimate) ? 237:
			/**/
			/**/
			 /**/
			(r_counter == 118 & r_state==zStateEstimate) ? 668:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 120 & r_state==zStateEstimate) ? 238:
			/**/
			/**/
			 /**/
			(r_counter == 121 & r_state==zStateEstimate) ? 497:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 123 & r_state==zStateEstimate) ? 121:
			/**/
			/**/
			 /**/
			(r_counter == 124 & r_state==zStateEstimate) ? 712:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 126 & r_state==zStateEstimate) ? 240:
			/**/
			/**/
			 /**/
			(r_counter == 127 & r_state==zStateEstimate) ? 696:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 129 & r_state==zStateEstimate) ? 241:
			/**/
			/**/
			 /**/
			(r_counter == 130 & r_state==zStateEstimate) ? 600:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 132 & r_state==zStateEstimate) ? 242:
			/**/
			/**/
			 /**/
			(r_counter == 133 & r_state==zStateEstimate) ? 764:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 135 & r_state==zStateEstimate) ? 156:
			/**/
			/**/
			 /**/
			(r_counter == 136 & r_state==zStateEstimate) ? 516:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 138 & r_state==zStateEstimate) ? 244:
			/**/
			/**/
			 /**/
			(r_counter == 139 & r_state==zStateEstimate) ? 428:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 141 & r_state==zStateEstimate) ? 245:
			/**/
			/**/
			 /**/
			(r_counter == 142 & r_state==zStateEstimate) ? 725:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 144 & r_state==zStateEstimate) ? 246:
			/**/
			/**/
			 /**/
			(r_counter == 145 & r_state==zStateEstimate) ? 576:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 147 & r_state==zStateEstimate) ? 122:
			/**/
			/**/
			 /**/
			(r_counter == 148 & r_state==zStateEstimate) ? 556:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 150 & r_state==zStateEstimate) ? 248:
			/**/
			/**/
			 /**/
			(r_counter == 151 & r_state==zStateEstimate) ? 492:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 153 & r_state==zStateEstimate) ? 249:
			/**/
			/**/
			 /**/
			(r_counter == 154 & r_state==zStateEstimate) ? 632:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 156 & r_state==zStateEstimate) ? 250:
			/**/
			/**/
			 /**/
			(r_counter == 157 & r_state==zStateEstimate) ? 432:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 159 & r_state==zStateEstimate) ? 96:
			/**/
			/**/
			 /**/
			(r_counter == 160 & r_state==zStateEstimate) ? 508:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 162 & r_state==zStateEstimate) ? 97:
			/**/
			/**/
			 /**/
			(r_counter == 163 & r_state==zStateEstimate) ? 660:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 165 & r_state==zStateEstimate) ? 252:
			/**/
			/**/
			 /**/
			(r_counter == 166 & r_state==zStateEstimate) ? 672:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 168 & r_state==zStateEstimate) ? 253:
			/**/
			/**/
			 /**/
			(r_counter == 169 & r_state==zStateEstimate) ? 768:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 171 & r_state==zStateEstimate) ? 124:
			/**/
			/**/
			 /**/
			(r_counter == 172 & r_state==zStateEstimate) ? 577:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 174 & r_state==zStateEstimate) ? 256:
			/**/
			/**/
			 /**/
			(r_counter == 175 & r_state==zStateEstimate) ? 752:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 177 & r_state==zStateEstimate) ? 257:
			/**/
			/**/
			 /**/
			(r_counter == 178 & r_state==zStateEstimate) ? 528:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 180 & r_state==zStateEstimate) ? 258:
			/**/
			/**/
			 /**/
			(r_counter == 181 & r_state==zStateEstimate) ? 728:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 183 & r_state==zStateEstimate) ? 64:
			/**/
			/**/
			 /**/
			(r_counter == 184 & r_state==zStateEstimate) ? 448:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 186 & r_state==zStateEstimate) ? 260:
			/**/
			/**/
			 /**/
			(r_counter == 187 & r_state==zStateEstimate) ? 608:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 189 & r_state==zStateEstimate) ? 261:
			/**/
			/**/
			 /**/
			(r_counter == 190 & r_state==zStateEstimate) ? 748:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 192 & r_state==zStateEstimate) ? 262:
			/**/
			/**/
			 /**/
			(r_counter == 193 & r_state==zStateEstimate) ? 456:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 195 & r_state==zStateEstimate) ? 108:
			/**/
			/**/
			 /**/
			(r_counter == 196 & r_state==zStateEstimate) ? 429:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 198 & r_state==zStateEstimate) ? 264:
			/**/
			/**/
			 /**/
			(r_counter == 199 & r_state==zStateEstimate) ? 753:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 201 & r_state==zStateEstimate) ? 265:
			/**/
			/**/
			 /**/
			(r_counter == 202 & r_state==zStateEstimate) ? 529:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 204 & r_state==zStateEstimate) ? 266:
			/**/
			/**/
			 /**/
			(r_counter == 205 & r_state==zStateEstimate) ? 665:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 207 & r_state==zStateEstimate) ? 128:
			/**/
			/**/
			 /**/
			(r_counter == 208 & r_state==zStateEstimate) ? 417:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 210 & r_state==zStateEstimate) ? 268:
			/**/
			/**/
			 /**/
			(r_counter == 211 & r_state==zStateEstimate) ? 625:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 213 & r_state==zStateEstimate) ? 269:
			/**/
			/**/
			 /**/
			(r_counter == 214 & r_state==zStateEstimate) ? 700:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 216 & r_state==zStateEstimate) ? 270:
			/**/
			/**/
			 /**/
			(r_counter == 217 & r_state==zStateEstimate) ? 513:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 219 & r_state==zStateEstimate) ? 164:
			/**/
			/**/
			 /**/
			(r_counter == 220 & r_state==zStateEstimate) ? 765:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 222 & r_state==zStateEstimate) ? 272:
			/**/
			/**/
			 /**/
			(r_counter == 223 & r_state==zStateEstimate) ? 400:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 225 & r_state==zStateEstimate) ? 273:
			/**/
			/**/
			 /**/
			(r_counter == 226 & r_state==zStateEstimate) ? 769:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 228 & r_state==zStateEstimate) ? 274:
			/**/
			/**/
			 /**/
			(r_counter == 229 & r_state==zStateEstimate) ? 548:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 231 & r_state==zStateEstimate) ? 165:
			/**/
			/**/
			 /**/
			(r_counter == 232 & r_state==zStateEstimate) ? 749:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 234 & r_state==zStateEstimate) ? 276:
			/**/
			/**/
			 /**/
			(r_counter == 235 & r_state==zStateEstimate) ? 524:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 237 & r_state==zStateEstimate) ? 277:
			/**/
			/**/
			 /**/
			(r_counter == 238 & r_state==zStateEstimate) ? 473:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 240 & r_state==zStateEstimate) ? 278:
			/**/
			/**/
			 /**/
			(r_counter == 241 & r_state==zStateEstimate) ? 612:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 243 & r_state==zStateEstimate) ? 166:
			/**/
			/**/
			 /**/
			(r_counter == 244 & r_state==zStateEstimate) ? 708:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 246 & r_state==zStateEstimate) ? 280:
			/**/
			/**/
			 /**/
			(r_counter == 247 & r_state==zStateEstimate) ? 409:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 249 & r_state==zStateEstimate) ? 281:
			/**/
			/**/
			 /**/
			(r_counter == 250 & r_state==zStateEstimate) ? 796:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 252 & r_state==zStateEstimate) ? 282:
			/**/
			/**/
			 /**/
			(r_counter == 253 & r_state==zStateEstimate) ? 640:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 255 & r_state==zStateEstimate) ? 129:
			/**/
			/**/
			 /**/
			(r_counter == 256 & r_state==zStateEstimate) ? 797:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 258 & r_state==zStateEstimate) ? 284:
			/**/
			/**/
			 /**/
			(r_counter == 259 & r_state==zStateEstimate) ? 498:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 261 & r_state==zStateEstimate) ? 285:
			/**/
			/**/
			 /**/
			(r_counter == 262 & r_state==zStateEstimate) ? 744:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 264 & r_state==zStateEstimate) ? 286:
			/**/
			/**/
			 /**/
			(r_counter == 265 & r_state==zStateEstimate) ? 449:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 267 & r_state==zStateEstimate) ? 168:
			/**/
			/**/
			 /**/
			(r_counter == 268 & r_state==zStateEstimate) ? 532:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 270 & r_state==zStateEstimate) ? 288:
			/**/
			/**/
			 /**/
			(r_counter == 271 & r_state==zStateEstimate) ? 777:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 273 & r_state==zStateEstimate) ? 169:
			/**/
			/**/
			 /**/
			(r_counter == 274 & r_state==zStateEstimate) ? 717:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 276 & r_state==zStateEstimate) ? 289:
			/**/
			/**/
			 /**/
			(r_counter == 277 & r_state==zStateEstimate) ? 621:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 279 & r_state==zStateEstimate) ? 170:
			/**/
			/**/
			 /**/
			(r_counter == 280 & r_state==zStateEstimate) ? 736:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 282 & r_state==zStateEstimate) ? 292:
			/**/
			/**/
			 /**/
			(r_counter == 283 & r_state==zStateEstimate) ? 680:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 285 & r_state==zStateEstimate) ? 293:
			/**/
			/**/
			 /**/
			(r_counter == 286 & r_state==zStateEstimate) ? 505:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 288 & r_state==zStateEstimate) ? 294:
			/**/
			/**/
			 /**/
			(r_counter == 289 & r_state==zStateEstimate) ? 480:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 291 & r_state==zStateEstimate) ? 130:
			/**/
			/**/
			 /**/
			(r_counter == 292 & r_state==zStateEstimate) ? 756:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 294 & r_state==zStateEstimate) ? 296:
			/**/
			/**/
			 /**/
			(r_counter == 295 & r_state==zStateEstimate) ? 444:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 297 & r_state==zStateEstimate) ? 297:
			/**/
			/**/
			 /**/
			(r_counter == 298 & r_state==zStateEstimate) ? 500:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 300 & r_state==zStateEstimate) ? 298:
			/**/
			/**/
			 /**/
			(r_counter == 301 & r_state==zStateEstimate) ? 745:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 303 & r_state==zStateEstimate) ? 84:
			/**/
			/**/
			 /**/
			(r_counter == 304 & r_state==zStateEstimate) ? 433:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 306 & r_state==zStateEstimate) ? 300:
			/**/
			/**/
			 /**/
			(r_counter == 307 & r_state==zStateEstimate) ? 457:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 309 & r_state==zStateEstimate) ? 301:
			/**/
			/**/
			 /**/
			(r_counter == 310 & r_state==zStateEstimate) ? 729:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 312 & r_state==zStateEstimate) ? 302:
			/**/
			/**/
			 /**/
			(r_counter == 313 & r_state==zStateEstimate) ? 673:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 315 & r_state==zStateEstimate) ? 132:
			/**/
			/**/
			 /**/
			(r_counter == 316 & r_state==zStateEstimate) ? 468:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 318 & r_state==zStateEstimate) ? 304:
			/**/
			/**/
			 /**/
			(r_counter == 319 & r_state==zStateEstimate) ? 648:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 321 & r_state==zStateEstimate) ? 305:
			/**/
			/**/
			 /**/
			(r_counter == 322 & r_state==zStateEstimate) ? 549:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 324 & r_state==zStateEstimate) ? 306:
			/**/
			/**/
			 /**/
			(r_counter == 325 & r_state==zStateEstimate) ? 533:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 327 & r_state==zStateEstimate) ? 172:
			/**/
			/**/
			 /**/
			(r_counter == 328 & r_state==zStateEstimate) ? 701:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 330 & r_state==zStateEstimate) ? 133:
			/**/
			/**/
			 /**/
			(r_counter == 331 & r_state==zStateEstimate) ? 437:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 333 & r_state==zStateEstimate) ? 308:
			/**/
			/**/
			 /**/
			(r_counter == 334 & r_state==zStateEstimate) ? 780:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 336 & r_state==zStateEstimate) ? 309:
			/**/
			/**/
			 /**/
			(r_counter == 337 & r_state==zStateEstimate) ? 445:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 339 & r_state==zStateEstimate) ? 176:
			/**/
			/**/
			 /**/
			(r_counter == 340 & r_state==zStateEstimate) ? 412:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 342 & r_state==zStateEstimate) ? 312:
			/**/
			/**/
			 /**/
			(r_counter == 343 & r_state==zStateEstimate) ? 718:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 345 & r_state==zStateEstimate) ? 313:
			/**/
			/**/
			 /**/
			(r_counter == 346 & r_state==zStateEstimate) ? 674:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 348 & r_state==zStateEstimate) ? 314:
			/**/
			/**/
			 /**/
			(r_counter == 349 & r_state==zStateEstimate) ? 580:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 351 & r_state==zStateEstimate) ? 177:
			/**/
			/**/
			 /**/
			(r_counter == 352 & r_state==zStateEstimate) ? 684:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 354 & r_state==zStateEstimate) ? 316:
			/**/
			/**/
			 /**/
			(r_counter == 355 & r_state==zStateEstimate) ? 544:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 357 & r_state==zStateEstimate) ? 317:
			/**/
			/**/
			 /**/
			(r_counter == 358 & r_state==zStateEstimate) ? 484:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 360 & r_state==zStateEstimate) ? 318:
			/**/
			/**/
			 /**/
			(r_counter == 361 & r_state==zStateEstimate) ? 628:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 363 & r_state==zStateEstimate) ? 134:
			/**/
			/**/
			 /**/
			(r_counter == 364 & r_state==zStateEstimate) ? 713:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 366 & r_state==zStateEstimate) ? 320:
			/**/
			/**/
			 /**/
			(r_counter == 367 & r_state==zStateEstimate) ? 609:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 369 & r_state==zStateEstimate) ? 321:
			/**/
			/**/
			 /**/
			(r_counter == 370 & r_state==zStateEstimate) ? 645:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 372 & r_state==zStateEstimate) ? 322:
			/**/
			/**/
			 /**/
			(r_counter == 373 & r_state==zStateEstimate) ? 692:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 375 & r_state==zStateEstimate) ? 0:
			/**/
			/**/
			 /**/
			(r_counter == 376 & r_state==zStateEstimate) ? 565:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 378 & r_state==zStateEstimate) ? 324:
			/**/
			/**/
			 /**/
			(r_counter == 379 & r_state==zStateEstimate) ? 413:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 381 & r_state==zStateEstimate) ? 325:
			/**/
			/**/
			 /**/
			(r_counter == 382 & r_state==zStateEstimate) ? 585:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 384 & r_state==zStateEstimate) ? 326:
			/**/
			/**/
			 /**/
			(r_counter == 385 & r_state==zStateEstimate) ? 661:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 387 & r_state==zStateEstimate) ? 136:
			/**/
			/**/
			 /**/
			(r_counter == 388 & r_state==zStateEstimate) ? 485:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 390 & r_state==zStateEstimate) ? 328:
			/**/
			/**/
			 /**/
			(r_counter == 391 & r_state==zStateEstimate) ? 450:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 393 & r_state==zStateEstimate) ? 329:
			/**/
			/**/
			 /**/
			(r_counter == 394 & r_state==zStateEstimate) ? 452:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 396 & r_state==zStateEstimate) ? 330:
			/**/
			/**/
			 /**/
			(r_counter == 397 & r_state==zStateEstimate) ? 633:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 399 & r_state==zStateEstimate) ? 137:
			/**/
			/**/
			 /**/
			(r_counter == 400 & r_state==zStateEstimate) ? 662:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 402 & r_state==zStateEstimate) ? 332:
			/**/
			/**/
			 /**/
			(r_counter == 403 & r_state==zStateEstimate) ? 720:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 405 & r_state==zStateEstimate) ? 333:
			/**/
			/**/
			 /**/
			(r_counter == 406 & r_state==zStateEstimate) ? 401:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 408 & r_state==zStateEstimate) ? 334:
			/**/
			/**/
			 /**/
			(r_counter == 409 & r_state==zStateEstimate) ? 481:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 411 & r_state==zStateEstimate) ? 180:
			/**/
			/**/
			 /**/
			(r_counter == 412 & r_state==zStateEstimate) ? 493:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 414 & r_state==zStateEstimate) ? 336:
			/**/
			/**/
			 /**/
			(r_counter == 415 & r_state==zStateEstimate) ? 634:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 417 & r_state==zStateEstimate) ? 337:
			/**/
			/**/
			 /**/
			(r_counter == 418 & r_state==zStateEstimate) ? 721:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 420 & r_state==zStateEstimate) ? 338:
			/**/
			/**/
			 /**/
			(r_counter == 421 & r_state==zStateEstimate) ? 568:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 423 & r_state==zStateEstimate) ? 138:
			/**/
			/**/
			 /**/
			(r_counter == 424 & r_state==zStateEstimate) ? 733:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 426 & r_state==zStateEstimate) ? 340:
			/**/
			/**/
			 /**/
			(r_counter == 427 & r_state==zStateEstimate) ? 588:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 429 & r_state==zStateEstimate) ? 341:
			/**/
			/**/
			 /**/
			(r_counter == 430 & r_state==zStateEstimate) ? 610:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 432 & r_state==zStateEstimate) ? 342:
			/**/
			/**/
			 /**/
			(r_counter == 433 & r_state==zStateEstimate) ? 545:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 435 & r_state==zStateEstimate) ? 184:
			/**/
			/**/
			 /**/
			(r_counter == 436 & r_state==zStateEstimate) ? 629:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 438 & r_state==zStateEstimate) ? 344:
			/**/
			/**/
			 /**/
			(r_counter == 439 & r_state==zStateEstimate) ? 569:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 441 & r_state==zStateEstimate) ? 345:
			/**/
			/**/
			 /**/
			(r_counter == 442 & r_state==zStateEstimate) ? 778:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 444 & r_state==zStateEstimate) ? 346:
			/**/
			/**/
			 /**/
			(r_counter == 445 & r_state==zStateEstimate) ? 754:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 447 & r_state==zStateEstimate) ? 185:
			/**/
			/**/
			 /**/
			(r_counter == 448 & r_state==zStateEstimate) ? 709:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 450 & r_state==zStateEstimate) ? 348:
			/**/
			/**/
			 /**/
			(r_counter == 451 & r_state==zStateEstimate) ? 477:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 453 & r_state==zStateEstimate) ? 349:
			/**/
			/**/
			 /**/
			(r_counter == 454 & r_state==zStateEstimate) ? 546:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 456 & r_state==zStateEstimate) ? 350:
			/**/
			/**/
			 /**/
			(r_counter == 457 & r_state==zStateEstimate) ? 586:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 459 & r_state==zStateEstimate) ? 186:
			/**/
			/**/
			 /**/
			(r_counter == 460 & r_state==zStateEstimate) ? 536:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 462 & r_state==zStateEstimate) ? 352:
			/**/
			/**/
			 /**/
			(r_counter == 463 & r_state==zStateEstimate) ? 613:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 465 & r_state==zStateEstimate) ? 353:
			/**/
			/**/
			 /**/
			(r_counter == 466 & r_state==zStateEstimate) ? 652:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 468 & r_state==zStateEstimate) ? 354:
			/**/
			/**/
			 /**/
			(r_counter == 469 & r_state==zStateEstimate) ? 622:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 471 & r_state==zStateEstimate) ? 100:
			/**/
			/**/
			 /**/
			(r_counter == 472 & r_state==zStateEstimate) ? 702:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 474 & r_state==zStateEstimate) ? 356:
			/**/
			/**/
			 /**/
			(r_counter == 475 & r_state==zStateEstimate) ? 592:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 477 & r_state==zStateEstimate) ? 357:
			/**/
			/**/
			 /**/
			(r_counter == 478 & r_state==zStateEstimate) ? 760:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 480 & r_state==zStateEstimate) ? 358:
			/**/
			/**/
			 /**/
			(r_counter == 481 & r_state==zStateEstimate) ? 630:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 483 & r_state==zStateEstimate) ? 188:
			/**/
			/**/
			 /**/
			(r_counter == 484 & r_state==zStateEstimate) ? 440:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 486 & r_state==zStateEstimate) ? 360:
			/**/
			/**/
			 /**/
			(r_counter == 487 & r_state==zStateEstimate) ? 557:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 489 & r_state==zStateEstimate) ? 361:
			/**/
			/**/
			 /**/
			(r_counter == 490 & r_state==zStateEstimate) ? 693:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 492 & r_state==zStateEstimate) ? 362:
			/**/
			/**/
			 /**/
			(r_counter == 493 & r_state==zStateEstimate) ? 637:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 495 & r_state==zStateEstimate) ? 189:
			/**/
			/**/
			 /**/
			(r_counter == 496 & r_state==zStateEstimate) ? 677:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 498 & r_state==zStateEstimate) ? 364:
			/**/
			/**/
			 /**/
			(r_counter == 499 & r_state==zStateEstimate) ? 596:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 501 & r_state==zStateEstimate) ? 365:
			/**/
			/**/
			 /**/
			(r_counter == 502 & r_state==zStateEstimate) ? 616:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 504 & r_state==zStateEstimate) ? 366:
			/**/
			/**/
			 /**/
			(r_counter == 505 & r_state==zStateEstimate) ? 520:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 507 & r_state==zStateEstimate) ? 190:
			/**/
			/**/
			 /**/
			(r_counter == 508 & r_state==zStateEstimate) ? 705:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 510 & r_state==zStateEstimate) ? 368:
			/**/
			/**/
			 /**/
			(r_counter == 511 & r_state==zStateEstimate) ? 578:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 513 & r_state==zStateEstimate) ? 369:
			/**/
			/**/
			 /**/
			(r_counter == 514 & r_state==zStateEstimate) ? 617:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 516 & r_state==zStateEstimate) ? 370:
			/**/
			/**/
			 /**/
			(r_counter == 517 & r_state==zStateEstimate) ? 641:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 519 & r_state==zStateEstimate) ? 113:
			/**/
			/**/
			 /**/
			(r_counter == 520 & r_state==zStateEstimate) ? 488:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 522 & r_state==zStateEstimate) ? 372:
			/**/
			/**/
			 /**/
			(r_counter == 523 & r_state==zStateEstimate) ? 446:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 525 & r_state==zStateEstimate) ? 373:
			/**/
			/**/
			 /**/
			(r_counter == 526 & r_state==zStateEstimate) ? 685:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 528 & r_state==zStateEstimate) ? 374:
			/**/
			/**/
			 /**/
			(r_counter == 529 & r_state==zStateEstimate) ? 741:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 531 & r_state==zStateEstimate) ? 192:
			/**/
			/**/
			 /**/
			(r_counter == 532 & r_state==zStateEstimate) ? 726:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 534 & r_state==zStateEstimate) ? 376:
			/**/
			/**/
			 /**/
			(r_counter == 535 & r_state==zStateEstimate) ? 402:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 537 & r_state==zStateEstimate) ? 377:
			/**/
			/**/
			 /**/
			(r_counter == 538 & r_state==zStateEstimate) ? 697:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 540 & r_state==zStateEstimate) ? 378:
			/**/
			/**/
			 /**/
			(r_counter == 541 & r_state==zStateEstimate) ? 466:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 543 & r_state==zStateEstimate) ? 193:
			/**/
			/**/
			 /**/
			(r_counter == 544 & r_state==zStateEstimate) ? 798:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 546 & r_state==zStateEstimate) ? 380:
			/**/
			/**/
			 /**/
			(r_counter == 547 & r_state==zStateEstimate) ? 521:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 549 & r_state==zStateEstimate) ? 381:
			/**/
			/**/
			 /**/
			(r_counter == 550 & r_state==zStateEstimate) ? 573:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 552 & r_state==zStateEstimate) ? 382:
			/**/
			/**/
			 /**/
			(r_counter == 553 & r_state==zStateEstimate) ? 506:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 555 & r_state==zStateEstimate) ? 194:
			/**/
			/**/
			 /**/
			(r_counter == 556 & r_state==zStateEstimate) ? 785:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 558 & r_state==zStateEstimate) ? 384:
			/**/
			/**/
			 /**/
			(r_counter == 559 & r_state==zStateEstimate) ? 781:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 561 & r_state==zStateEstimate) ? 385:
			/**/
			/**/
			 /**/
			(r_counter == 562 & r_state==zStateEstimate) ? 530:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 564 & r_state==zStateEstimate) ? 386:
			/**/
			/**/
			 /**/
			(r_counter == 565 & r_state==zStateEstimate) ? 589:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 567 & r_state==zStateEstimate) ? 141:
			/**/
			/**/
			 /**/
			(r_counter == 568 & r_state==zStateEstimate) ? 424:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 570 & r_state==zStateEstimate) ? 388:
			/**/
			/**/
			 /**/
			(r_counter == 571 & r_state==zStateEstimate) ? 525:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 573 & r_state==zStateEstimate) ? 389:
			/**/
			/**/
			 /**/
			(r_counter == 574 & r_state==zStateEstimate) ? 761:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 576 & r_state==zStateEstimate) ? 390:
			/**/
			/**/
			 /**/
			(r_counter == 577 & r_state==zStateEstimate) ? 618:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 579 & r_state==zStateEstimate) ? 197:
			/**/
			/**/
			 /**/
			(r_counter == 580 & r_state==zStateEstimate) ? 793:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 582 & r_state==zStateEstimate) ? 392:
			/**/
			/**/
			 /**/
			(r_counter == 583 & r_state==zStateEstimate) ? 478:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 585 & r_state==zStateEstimate) ? 393:
			/**/
			/**/
			 /**/
			(r_counter == 586 & r_state==zStateEstimate) ? 482:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 588 & r_state==zStateEstimate) ? 394:
			/**/
			/**/
			 /**/
			(r_counter == 589 & r_state==zStateEstimate) ? 438:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 591 & r_state==zStateEstimate) ? 198:
			/**/
			/**/
			 /**/
			(r_counter == 592 & r_state==zStateEstimate) ? 601:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 594 & r_state==zStateEstimate) ? 396:
			/**/
			/**/
			 /**/
			(r_counter == 595 & r_state==zStateEstimate) ? 421:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 597 & r_state==zStateEstimate) ? 397:
			/**/
			/**/
			 /**/
			(r_counter == 598 & r_state==zStateEstimate) ? 453:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 600 & r_state==zStateEstimate) ? 398:
			/**/
			/**/
			 /**/
			(r_counter == 601 & r_state==zStateEstimate) ? 653:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 603 & r_state==zStateEstimate) ? 1:
			/**/
			/**/
			 /**/
			(r_counter == 604 & r_state==zStateEstimate) ? 566:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 606 & r_state==zStateEstimate) ? 2:
			/**/
			/**/
			 /**/
			(r_counter == 607 & r_state==zStateEstimate) ? 489:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 609 & r_state==zStateEstimate) ? 3:
			/**/
			/**/
			 /**/
			(r_counter == 610 & r_state==zStateEstimate) ? 678:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 612 & r_state==zStateEstimate) ? 4:
			/**/
			/**/
			 /**/
			(r_counter == 613 & r_state==zStateEstimate) ? 794:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 615 & r_state==zStateEstimate) ? 5:
			/**/
			/**/
			 /**/
			(r_counter == 616 & r_state==zStateEstimate) ? 404:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 618 & r_state==zStateEstimate) ? 6:
			/**/
			/**/
			 /**/
			(r_counter == 619 & r_state==zStateEstimate) ? 509:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 621 & r_state==zStateEstimate) ? 7:
			/**/
			/**/
			 /**/
			(r_counter == 622 & r_state==zStateEstimate) ? 422:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 624 & r_state==zStateEstimate) ? 8:
			/**/
			/**/
			 /**/
			(r_counter == 625 & r_state==zStateEstimate) ? 642:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 627 & r_state==zStateEstimate) ? 9:
			/**/
			/**/
			 /**/
			(r_counter == 628 & r_state==zStateEstimate) ? 561:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 630 & r_state==zStateEstimate) ? 10:
			/**/
			/**/
			 /**/
			(r_counter == 631 & r_state==zStateEstimate) ? 434:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 633 & r_state==zStateEstimate) ? 11:
			/**/
			/**/
			 /**/
			(r_counter == 634 & r_state==zStateEstimate) ? 657:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 636 & r_state==zStateEstimate) ? 12:
			/**/
			/**/
			 /**/
			(r_counter == 637 & r_state==zStateEstimate) ? 517:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 639 & r_state==zStateEstimate) ? 13:
			/**/
			/**/
			 /**/
			(r_counter == 640 & r_state==zStateEstimate) ? 537:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 642 & r_state==zStateEstimate) ? 14:
			/**/
			/**/
			 /**/
			(r_counter == 643 & r_state==zStateEstimate) ? 554:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 645 & r_state==zStateEstimate) ? 15:
			/**/
			/**/
			 /**/
			(r_counter == 646 & r_state==zStateEstimate) ? 766:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 648 & r_state==zStateEstimate) ? 16:
			/**/
			/**/
			 /**/
			(r_counter == 649 & r_state==zStateEstimate) ? 719:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 651 & r_state==zStateEstimate) ? 17:
			/**/
			/**/
			 /**/
			(r_counter == 652 & r_state==zStateEstimate) ? 646:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 654 & r_state==zStateEstimate) ? 18:
			/**/
			/**/
			 /**/
			(r_counter == 655 & r_state==zStateEstimate) ? 593:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 657 & r_state==zStateEstimate) ? 19:
			/**/
			/**/
			 /**/
			(r_counter == 658 & r_state==zStateEstimate) ? 602:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 660 & r_state==zStateEstimate) ? 20:
			/**/
			/**/
			 /**/
			(r_counter == 661 & r_state==zStateEstimate) ? 666:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 663 & r_state==zStateEstimate) ? 21:
			/**/
			/**/
			 /**/
			(r_counter == 664 & r_state==zStateEstimate) ? 501:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 666 & r_state==zStateEstimate) ? 22:
			/**/
			/**/
			 /**/
			(r_counter == 667 & r_state==zStateEstimate) ? 737:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 669 & r_state==zStateEstimate) ? 23:
			/**/
			/**/
			 /**/
			(r_counter == 670 & r_state==zStateEstimate) ? 490:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 672 & r_state==zStateEstimate) ? 24:
			/**/
			/**/
			 /**/
			(r_counter == 673 & r_state==zStateEstimate) ? 558:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 675 & r_state==zStateEstimate) ? 25:
			/**/
			/**/
			 /**/
			(r_counter == 676 & r_state==zStateEstimate) ? 706:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 678 & r_state==zStateEstimate) ? 26:
			/**/
			/**/
			 /**/
			(r_counter == 679 & r_state==zStateEstimate) ? 474:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 681 & r_state==zStateEstimate) ? 27:
			/**/
			/**/
			 /**/
			(r_counter == 682 & r_state==zStateEstimate) ? 635:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 684 & r_state==zStateEstimate) ? 28:
			/**/
			/**/
			 /**/
			(r_counter == 685 & r_state==zStateEstimate) ? 469:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 687 & r_state==zStateEstimate) ? 29:
			/**/
			/**/
			 /**/
			(r_counter == 688 & r_state==zStateEstimate) ? 494:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 690 & r_state==zStateEstimate) ? 30:
			/**/
			/**/
			 /**/
			(r_counter == 691 & r_state==zStateEstimate) ? 714:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 693 & r_state==zStateEstimate) ? 31:
			/**/
			/**/
			 /**/
			(r_counter == 694 & r_state==zStateEstimate) ? 605:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 696 & r_state==zStateEstimate) ? 32:
			/**/
			/**/
			 /**/
			(r_counter == 697 & r_state==zStateEstimate) ? 707:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 699 & r_state==zStateEstimate) ? 33:
			/**/
			/**/
			 /**/
			(r_counter == 700 & r_state==zStateEstimate) ? 643:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 702 & r_state==zStateEstimate) ? 34:
			/**/
			/**/
			 /**/
			(r_counter == 703 & r_state==zStateEstimate) ? 579:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 705 & r_state==zStateEstimate) ? 35:
			/**/
			/**/
			 /**/
			(r_counter == 706 & r_state==zStateEstimate) ? 770:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 708 & r_state==zStateEstimate) ? 36:
			/**/
			/**/
			 /**/
			(r_counter == 709 & r_state==zStateEstimate) ? 405:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 711 & r_state==zStateEstimate) ? 37:
			/**/
			/**/
			 /**/
			(r_counter == 712 & r_state==zStateEstimate) ? 779:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 714 & r_state==zStateEstimate) ? 38:
			/**/
			/**/
			 /**/
			(r_counter == 715 & r_state==zStateEstimate) ? 514:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 717 & r_state==zStateEstimate) ? 39:
			/**/
			/**/
			 /**/
			(r_counter == 718 & r_state==zStateEstimate) ? 581:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 720 & r_state==zStateEstimate) ? 40:
			/**/
			/**/
			 /**/
			(r_counter == 721 & r_state==zStateEstimate) ? 746:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 723 & r_state==zStateEstimate) ? 41:
			/**/
			/**/
			 /**/
			(r_counter == 724 & r_state==zStateEstimate) ? 611:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 726 & r_state==zStateEstimate) ? 42:
			/**/
			/**/
			 /**/
			(r_counter == 727 & r_state==zStateEstimate) ? 510:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 729 & r_state==zStateEstimate) ? 43:
			/**/
			/**/
			 /**/
			(r_counter == 730 & r_state==zStateEstimate) ? 467:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 732 & r_state==zStateEstimate) ? 44:
			/**/
			/**/
			 /**/
			(r_counter == 733 & r_state==zStateEstimate) ? 502:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 735 & r_state==zStateEstimate) ? 45:
			/**/
			/**/
			 /**/
			(r_counter == 736 & r_state==zStateEstimate) ? 742:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 738 & r_state==zStateEstimate) ? 46:
			/**/
			/**/
			 /**/
			(r_counter == 739 & r_state==zStateEstimate) ? 538:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 741 & r_state==zStateEstimate) ? 47:
			/**/
			/**/
			 /**/
			(r_counter == 742 & r_state==zStateEstimate) ? 786:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 744 & r_state==zStateEstimate) ? 49:
			/**/
			/**/
			 /**/
			(r_counter == 745 & r_state==zStateEstimate) ? 511:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 747 & r_state==zStateEstimate) ? 50:
			/**/
			/**/
			 /**/
			(r_counter == 748 & r_state==zStateEstimate) ? 597:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 750 & r_state==zStateEstimate) ? 51:
			/**/
			/**/
			 /**/
			(r_counter == 751 & r_state==zStateEstimate) ? 451:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 753 & r_state==zStateEstimate) ? 52:
			/**/
			/**/
			 /**/
			(r_counter == 754 & r_state==zStateEstimate) ? 518:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 756 & r_state==zStateEstimate) ? 53:
			/**/
			/**/
			 /**/
			(r_counter == 757 & r_state==zStateEstimate) ? 486:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 759 & r_state==zStateEstimate) ? 54:
			/**/
			/**/
			 /**/
			(r_counter == 760 & r_state==zStateEstimate) ? 734:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 762 & r_state==zStateEstimate) ? 55:
			/**/
			/**/
			 /**/
			(r_counter == 763 & r_state==zStateEstimate) ? 460:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 765 & r_state==zStateEstimate) ? 56:
			/**/
			/**/
			 /**/
			(r_counter == 766 & r_state==zStateEstimate) ? 690:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 768 & r_state==zStateEstimate) ? 57:
			/**/
			/**/
			 /**/
			(r_counter == 769 & r_state==zStateEstimate) ? 799:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 771 & r_state==zStateEstimate) ? 58:
			/**/
			/**/
			 /**/
			(r_counter == 772 & r_state==zStateEstimate) ? 439:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 774 & r_state==zStateEstimate) ? 59:
			/**/
			/**/
			 /**/
			(r_counter == 775 & r_state==zStateEstimate) ? 425:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 777 & r_state==zStateEstimate) ? 60:
			/**/
			/**/
			 /**/
			(r_counter == 778 & r_state==zStateEstimate) ? 727:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 780 & r_state==zStateEstimate) ? 61:
			/**/
			/**/
			 /**/
			(r_counter == 781 & r_state==zStateEstimate) ? 638:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 783 & r_state==zStateEstimate) ? 62:
			/**/
			/**/
			 /**/
			(r_counter == 784 & r_state==zStateEstimate) ? 541:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 786 & r_state==zStateEstimate) ? 63:
			/**/
			/**/
			 /**/
			(r_counter == 787 & r_state==zStateEstimate) ? 658:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 789 & r_state==zStateEstimate) ? 65:
			/**/
			/**/
			 /**/
			(r_counter == 790 & r_state==zStateEstimate) ? 675:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 792 & r_state==zStateEstimate) ? 66:
			/**/
			/**/
			 /**/
			(r_counter == 793 & r_state==zStateEstimate) ? 774:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 795 & r_state==zStateEstimate) ? 67:
			/**/
			/**/
			 /**/
			(r_counter == 796 & r_state==zStateEstimate) ? 747:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 798 & r_state==zStateEstimate) ? 68:
			/**/
			/**/
			 /**/
			(r_counter == 799 & r_state==zStateEstimate) ? 594:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 801 & r_state==zStateEstimate) ? 69:
			/**/
			/**/
			 /**/
			(r_counter == 802 & r_state==zStateEstimate) ? 503:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 804 & r_state==zStateEstimate) ? 70:
			/**/
			/**/
			 /**/
			(r_counter == 805 & r_state==zStateEstimate) ? 694:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 807 & r_state==zStateEstimate) ? 71:
			/**/
			/**/
			 /**/
			(r_counter == 808 & r_state==zStateEstimate) ? 663:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 810 & r_state==zStateEstimate) ? 73:
			/**/
			/**/
			 /**/
			(r_counter == 811 & r_state==zStateEstimate) ? 542:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 813 & r_state==zStateEstimate) ? 74:
			/**/
			/**/
			 /**/
			(r_counter == 814 & r_state==zStateEstimate) ? 426:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 816 & r_state==zStateEstimate) ? 75:
			/**/
			/**/
			 /**/
			(r_counter == 817 & r_state==zStateEstimate) ? 495:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 819 & r_state==zStateEstimate) ? 76:
			/**/
			/**/
			 /**/
			(r_counter == 820 & r_state==zStateEstimate) ? 562:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 822 & r_state==zStateEstimate) ? 77:
			/**/
			/**/
			 /**/
			(r_counter == 823 & r_state==zStateEstimate) ? 534:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 825 & r_state==zStateEstimate) ? 78:
			/**/
			/**/
			 /**/
			(r_counter == 826 & r_state==zStateEstimate) ? 619:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 828 & r_state==zStateEstimate) ? 79:
			/**/
			/**/
			 /**/
			(r_counter == 829 & r_state==zStateEstimate) ? 598:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 831 & r_state==zStateEstimate) ? 80:
			/**/
			/**/
			 /**/
			(r_counter == 832 & r_state==zStateEstimate) ? 441:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 834 & r_state==zStateEstimate) ? 81:
			/**/
			/**/
			 /**/
			(r_counter == 835 & r_state==zStateEstimate) ? 606:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 837 & r_state==zStateEstimate) ? 82:
			/**/
			/**/
			 /**/
			(r_counter == 838 & r_state==zStateEstimate) ? 669:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 840 & r_state==zStateEstimate) ? 83:
			/**/
			/**/
			 /**/
			(r_counter == 841 & r_state==zStateEstimate) ? 479:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 843 & r_state==zStateEstimate) ? 85:
			/**/
			/**/
			 /**/
			(r_counter == 844 & r_state==zStateEstimate) ? 750:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 846 & r_state==zStateEstimate) ? 86:
			/**/
			/**/
			 /**/
			(r_counter == 847 & r_state==zStateEstimate) ? 735:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 849 & r_state==zStateEstimate) ? 87:
			/**/
			/**/
			 /**/
			(r_counter == 850 & r_state==zStateEstimate) ? 543:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 852 & r_state==zStateEstimate) ? 89:
			/**/
			/**/
			 /**/
			(r_counter == 853 & r_state==zStateEstimate) ? 703:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 855 & r_state==zStateEstimate) ? 90:
			/**/
			/**/
			 /**/
			(r_counter == 856 & r_state==zStateEstimate) ? 406:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 858 & r_state==zStateEstimate) ? 91:
			/**/
			/**/
			 /**/
			(r_counter == 859 & r_state==zStateEstimate) ? 526:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 861 & r_state==zStateEstimate) ? 92:
			/**/
			/**/
			 /**/
			(r_counter == 862 & r_state==zStateEstimate) ? 698:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 864 & r_state==zStateEstimate) ? 93:
			/**/
			/**/
			 /**/
			(r_counter == 865 & r_state==zStateEstimate) ? 654:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 867 & r_state==zStateEstimate) ? 94:
			/**/
			/**/
			 /**/
			(r_counter == 868 & r_state==zStateEstimate) ? 710:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 870 & r_state==zStateEstimate) ? 95:
			/**/
			/**/
			 /**/
			(r_counter == 871 & r_state==zStateEstimate) ? 603:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 873 & r_state==zStateEstimate) ? 98:
			/**/
			/**/
			 /**/
			(r_counter == 874 & r_state==zStateEstimate) ? 639:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 876 & r_state==zStateEstimate) ? 99:
			/**/
			/**/
			 /**/
			(r_counter == 877 & r_state==zStateEstimate) ? 550:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 879 & r_state==zStateEstimate) ? 101:
			/**/
			/**/
			 /**/
			(r_counter == 880 & r_state==zStateEstimate) ? 499:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 882 & r_state==zStateEstimate) ? 102:
			/**/
			/**/
			 /**/
			(r_counter == 883 & r_state==zStateEstimate) ? 555:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 885 & r_state==zStateEstimate) ? 103:
			/**/
			/**/
			 /**/
			(r_counter == 886 & r_state==zStateEstimate) ? 418:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 888 & r_state==zStateEstimate) ? 104:
			/**/
			/**/
			 /**/
			(r_counter == 889 & r_state==zStateEstimate) ? 475:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 891 & r_state==zStateEstimate) ? 105:
			/**/
			/**/
			 /**/
			(r_counter == 892 & r_state==zStateEstimate) ? 649:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 894 & r_state==zStateEstimate) ? 106:
			/**/
			/**/
			 /**/
			(r_counter == 895 & r_state==zStateEstimate) ? 414:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 897 & r_state==zStateEstimate) ? 107:
			/**/
			/**/
			 /**/
			(r_counter == 898 & r_state==zStateEstimate) ? 522:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 900 & r_state==zStateEstimate) ? 109:
			/**/
			/**/
			 /**/
			(r_counter == 901 & r_state==zStateEstimate) ? 430:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 903 & r_state==zStateEstimate) ? 110:
			/**/
			/**/
			 /**/
			(r_counter == 904 & r_state==zStateEstimate) ? 626:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 906 & r_state==zStateEstimate) ? 111:
			/**/
			/**/
			 /**/
			(r_counter == 907 & r_state==zStateEstimate) ? 679:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 909 & r_state==zStateEstimate) ? 114:
			/**/
			/**/
			 /**/
			(r_counter == 910 & r_state==zStateEstimate) ? 647:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 912 & r_state==zStateEstimate) ? 115:
			/**/
			/**/
			 /**/
			(r_counter == 913 & r_state==zStateEstimate) ? 789:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 915 & r_state==zStateEstimate) ? 118:
			/**/
			/**/
			 /**/
			(r_counter == 916 & r_state==zStateEstimate) ? 715:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 918 & r_state==zStateEstimate) ? 119:
			/**/
			/**/
			 /**/
			(r_counter == 919 & r_state==zStateEstimate) ? 755:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 921 & r_state==zStateEstimate) ? 123:
			/**/
			/**/
			 /**/
			(r_counter == 922 & r_state==zStateEstimate) ? 771:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 924 & r_state==zStateEstimate) ? 125:
			/**/
			/**/
			 /**/
			(r_counter == 925 & r_state==zStateEstimate) ? 757:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 927 & r_state==zStateEstimate) ? 126:
			/**/
			/**/
			 /**/
			(r_counter == 928 & r_state==zStateEstimate) ? 767:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 930 & r_state==zStateEstimate) ? 127:
			/**/
			/**/
			 /**/
			(r_counter == 931 & r_state==zStateEstimate) ? 574:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 933 & r_state==zStateEstimate) ? 131:
			/**/
			/**/
			 /**/
			(r_counter == 934 & r_state==zStateEstimate) ? 795:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 936 & r_state==zStateEstimate) ? 135:
			/**/
			/**/
			 /**/
			(r_counter == 937 & r_state==zStateEstimate) ? 442:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 939 & r_state==zStateEstimate) ? 139:
			/**/
			/**/
			 /**/
			(r_counter == 940 & r_state==zStateEstimate) ? 738:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 942 & r_state==zStateEstimate) ? 142:
			/**/
			/**/
			 /**/
			(r_counter == 943 & r_state==zStateEstimate) ? 627:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 945 & r_state==zStateEstimate) ? 143:
			/**/
			/**/
			 /**/
			(r_counter == 946 & r_state==zStateEstimate) ? 483:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 948 & r_state==zStateEstimate) ? 145:
			/**/
			/**/
			 /**/
			(r_counter == 949 & r_state==zStateEstimate) ? 739:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 951 & r_state==zStateEstimate) ? 146:
			/**/
			/**/
			 /**/
			(r_counter == 952 & r_state==zStateEstimate) ? 447:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 954 & r_state==zStateEstimate) ? 147:
			/**/
			/**/
			 /**/
			(r_counter == 955 & r_state==zStateEstimate) ? 730:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 957 & r_state==zStateEstimate) ? 150:
			/**/
			/**/
			 /**/
			(r_counter == 958 & r_state==zStateEstimate) ? 567:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 960 & r_state==zStateEstimate) ? 151:
			/**/
			/**/
			 /**/
			(r_counter == 961 & r_state==zStateEstimate) ? 570:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 963 & r_state==zStateEstimate) ? 154:
			/**/
			/**/
			 /**/
			(r_counter == 964 & r_state==zStateEstimate) ? 699:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 966 & r_state==zStateEstimate) ? 155:
			/**/
			/**/
			 /**/
			(r_counter == 967 & r_state==zStateEstimate) ? 686:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 969 & r_state==zStateEstimate) ? 157:
			/**/
			/**/
			 /**/
			(r_counter == 970 & r_state==zStateEstimate) ? 599:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 972 & r_state==zStateEstimate) ? 158:
			/**/
			/**/
			 /**/
			(r_counter == 973 & r_state==zStateEstimate) ? 458:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 975 & r_state==zStateEstimate) ? 159:
			/**/
			/**/
			 /**/
			(r_counter == 976 & r_state==zStateEstimate) ? 403:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 978 & r_state==zStateEstimate) ? 160:
			/**/
			/**/
			 /**/
			(r_counter == 979 & r_state==zStateEstimate) ? 614:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 981 & r_state==zStateEstimate) ? 161:
			/**/
			/**/
			 /**/
			(r_counter == 982 & r_state==zStateEstimate) ? 507:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 984 & r_state==zStateEstimate) ? 162:
			/**/
			/**/
			 /**/
			(r_counter == 985 & r_state==zStateEstimate) ? 587:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 987 & r_state==zStateEstimate) ? 163:
			/**/
			/**/
			 /**/
			(r_counter == 988 & r_state==zStateEstimate) ? 415:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 990 & r_state==zStateEstimate) ? 167:
			/**/
			/**/
			 /**/
			(r_counter == 991 & r_state==zStateEstimate) ? 551:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 993 & r_state==zStateEstimate) ? 171:
			/**/
			/**/
			 /**/
			(r_counter == 994 & r_state==zStateEstimate) ? 470:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 996 & r_state==zStateEstimate) ? 173:
			/**/
			/**/
			 /**/
			(r_counter == 997 & r_state==zStateEstimate) ? 423:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 999 & r_state==zStateEstimate) ? 174:
			/**/
			/**/
			 /**/
			(r_counter == 1000 & r_state==zStateEstimate) ? 722:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1002 & r_state==zStateEstimate) ? 175:
			/**/
			/**/
			 /**/
			(r_counter == 1003 & r_state==zStateEstimate) ? 410:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1005 & r_state==zStateEstimate) ? 178:
			/**/
			/**/
			 /**/
			(r_counter == 1006 & r_state==zStateEstimate) ? 407:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1008 & r_state==zStateEstimate) ? 179:
			/**/
			/**/
			 /**/
			(r_counter == 1009 & r_state==zStateEstimate) ? 762:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1011 & r_state==zStateEstimate) ? 181:
			/**/
			/**/
			 /**/
			(r_counter == 1012 & r_state==zStateEstimate) ? 631:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1014 & r_state==zStateEstimate) ? 182:
			/**/
			/**/
			 /**/
			(r_counter == 1015 & r_state==zStateEstimate) ? 731:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1017 & r_state==zStateEstimate) ? 183:
			/**/
			/**/
			 /**/
			(r_counter == 1018 & r_state==zStateEstimate) ? 623:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1020 & r_state==zStateEstimate) ? 187:
			/**/
			/**/
			 /**/
			(r_counter == 1021 & r_state==zStateEstimate) ? 787:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1023 & r_state==zStateEstimate) ? 191:
			/**/
			/**/
			 /**/
			(r_counter == 1024 & r_state==zStateEstimate) ? 650:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1026 & r_state==zStateEstimate) ? 195:
			/**/
			/**/
			 /**/
			(r_counter == 1027 & r_state==zStateEstimate) ? 758:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1029 & r_state==zStateEstimate) ? 199:
			/**/
			/**/
			 /**/
			(r_counter == 1030 & r_state==zStateEstimate) ? 461:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1032 & r_state==zStateEstimate) ? 203:
			/**/
			/**/
			 /**/
			(r_counter == 1033 & r_state==zStateEstimate) ? 563:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1035 & r_state==zStateEstimate) ? 207:
			/**/
			/**/
			 /**/
			(r_counter == 1036 & r_state==zStateEstimate) ? 763:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1038 & r_state==zStateEstimate) ? 211:
			/**/
			/**/
			 /**/
			(r_counter == 1039 & r_state==zStateEstimate) ? 427:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1041 & r_state==zStateEstimate) ? 214:
			/**/
			/**/
			 /**/
			(r_counter == 1042 & r_state==zStateEstimate) ? 431:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1044 & r_state==zStateEstimate) ? 215:
			/**/
			/**/
			 /**/
			(r_counter == 1045 & r_state==zStateEstimate) ? 681:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1047 & r_state==zStateEstimate) ? 219:
			/**/
			/**/
			 /**/
			(r_counter == 1048 & r_state==zStateEstimate) ? 751:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1050 & r_state==zStateEstimate) ? 222:
			/**/
			/**/
			 /**/
			(r_counter == 1051 & r_state==zStateEstimate) ? 582:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1053 & r_state==zStateEstimate) ? 223:
			/**/
			/**/
			 /**/
			(r_counter == 1054 & r_state==zStateEstimate) ? 782:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1056 & r_state==zStateEstimate) ? 227:
			/**/
			/**/
			 /**/
			(r_counter == 1057 & r_state==zStateEstimate) ? 595:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1059 & r_state==zStateEstimate) ? 230:
			/**/
			/**/
			 /**/
			(r_counter == 1060 & r_state==zStateEstimate) ? 487:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1062 & r_state==zStateEstimate) ? 231:
			/**/
			/**/
			 /**/
			(r_counter == 1063 & r_state==zStateEstimate) ? 531:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1065 & r_state==zStateEstimate) ? 235:
			/**/
			/**/
			 /**/
			(r_counter == 1066 & r_state==zStateEstimate) ? 759:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1068 & r_state==zStateEstimate) ? 239:
			/**/
			/**/
			 /**/
			(r_counter == 1069 & r_state==zStateEstimate) ? 443:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1071 & r_state==zStateEstimate) ? 243:
			/**/
			/**/
			 /**/
			(r_counter == 1072 & r_state==zStateEstimate) ? 723:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1074 & r_state==zStateEstimate) ? 247:
			/**/
			/**/
			 /**/
			(r_counter == 1075 & r_state==zStateEstimate) ? 670:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1077 & r_state==zStateEstimate) ? 251:
			/**/
			/**/
			 /**/
			(r_counter == 1078 & r_state==zStateEstimate) ? 462:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1080 & r_state==zStateEstimate) ? 254:
			/**/
			/**/
			 /**/
			(r_counter == 1081 & r_state==zStateEstimate) ? 590:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1083 & r_state==zStateEstimate) ? 255:
			/**/
			/**/
			 /**/
			(r_counter == 1084 & r_state==zStateEstimate) ? 790:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1086 & r_state==zStateEstimate) ? 259:
			/**/
			/**/
			 /**/
			(r_counter == 1087 & r_state==zStateEstimate) ? 667:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1089 & r_state==zStateEstimate) ? 263:
			/**/
			/**/
			 /**/
			(r_counter == 1090 & r_state==zStateEstimate) ? 655:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1092 & r_state==zStateEstimate) ? 267:
			/**/
			/**/
			 /**/
			(r_counter == 1093 & r_state==zStateEstimate) ? 583:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1095 & r_state==zStateEstimate) ? 271:
			/**/
			/**/
			 /**/
			(r_counter == 1096 & r_state==zStateEstimate) ? 471:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1098 & r_state==zStateEstimate) ? 275:
			/**/
			/**/
			 /**/
			(r_counter == 1099 & r_state==zStateEstimate) ? 691:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1101 & r_state==zStateEstimate) ? 279:
			/**/
			/**/
			 /**/
			(r_counter == 1102 & r_state==zStateEstimate) ? 671:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1104 & r_state==zStateEstimate) ? 283:
			/**/
			/**/
			 /**/
			(r_counter == 1105 & r_state==zStateEstimate) ? 459:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1107 & r_state==zStateEstimate) ? 287:
			/**/
			/**/
			 /**/
			(r_counter == 1108 & r_state==zStateEstimate) ? 783:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1110 & r_state==zStateEstimate) ? 290:
			/**/
			/**/
			 /**/
			(r_counter == 1111 & r_state==zStateEstimate) ? 743:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1113 & r_state==zStateEstimate) ? 291:
			/**/
			/**/
			 /**/
			(r_counter == 1114 & r_state==zStateEstimate) ? 547:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1116 & r_state==zStateEstimate) ? 295:
			/**/
			/**/
			 /**/
			(r_counter == 1117 & r_state==zStateEstimate) ? 463:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1119 & r_state==zStateEstimate) ? 299:
			/**/
			/**/
			 /**/
			(r_counter == 1120 & r_state==zStateEstimate) ? 575:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1122 & r_state==zStateEstimate) ? 303:
			/**/
			/**/
			 /**/
			(r_counter == 1123 & r_state==zStateEstimate) ? 711:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1125 & r_state==zStateEstimate) ? 307:
			/**/
			/**/
			 /**/
			(r_counter == 1126 & r_state==zStateEstimate) ? 535:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1128 & r_state==zStateEstimate) ? 310:
			/**/
			/**/
			 /**/
			(r_counter == 1129 & r_state==zStateEstimate) ? 435:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1131 & r_state==zStateEstimate) ? 311:
			/**/
			/**/
			 /**/
			(r_counter == 1132 & r_state==zStateEstimate) ? 454:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1134 & r_state==zStateEstimate) ? 315:
			/**/
			/**/
			 /**/
			(r_counter == 1135 & r_state==zStateEstimate) ? 659:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1137 & r_state==zStateEstimate) ? 319:
			/**/
			/**/
			 /**/
			(r_counter == 1138 & r_state==zStateEstimate) ? 519:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1140 & r_state==zStateEstimate) ? 323:
			/**/
			/**/
			 /**/
			(r_counter == 1141 & r_state==zStateEstimate) ? 791:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1143 & r_state==zStateEstimate) ? 327:
			/**/
			/**/
			 /**/
			(r_counter == 1144 & r_state==zStateEstimate) ? 687:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1146 & r_state==zStateEstimate) ? 331:
			/**/
			/**/
			 /**/
			(r_counter == 1147 & r_state==zStateEstimate) ? 559:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1149 & r_state==zStateEstimate) ? 335:
			/**/
			/**/
			 /**/
			(r_counter == 1150 & r_state==zStateEstimate) ? 515:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1152 & r_state==zStateEstimate) ? 339:
			/**/
			/**/
			 /**/
			(r_counter == 1153 & r_state==zStateEstimate) ? 527:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1155 & r_state==zStateEstimate) ? 343:
			/**/
			/**/
			 /**/
			(r_counter == 1156 & r_state==zStateEstimate) ? 419:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1158 & r_state==zStateEstimate) ? 347:
			/**/
			/**/
			 /**/
			(r_counter == 1159 & r_state==zStateEstimate) ? 775:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1161 & r_state==zStateEstimate) ? 351:
			/**/
			/**/
			 /**/
			(r_counter == 1162 & r_state==zStateEstimate) ? 607:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1164 & r_state==zStateEstimate) ? 355:
			/**/
			/**/
			 /**/
			(r_counter == 1165 & r_state==zStateEstimate) ? 571:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1167 & r_state==zStateEstimate) ? 359:
			/**/
			/**/
			 /**/
			(r_counter == 1168 & r_state==zStateEstimate) ? 491:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1170 & r_state==zStateEstimate) ? 363:
			/**/
			/**/
			 /**/
			(r_counter == 1171 & r_state==zStateEstimate) ? 695:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1173 & r_state==zStateEstimate) ? 367:
			/**/
			/**/
			 /**/
			(r_counter == 1174 & r_state==zStateEstimate) ? 411:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1176 & r_state==zStateEstimate) ? 371:
			/**/
			/**/
			 /**/
			(r_counter == 1177 & r_state==zStateEstimate) ? 523:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1179 & r_state==zStateEstimate) ? 375:
			/**/
			/**/
			 /**/
			(r_counter == 1180 & r_state==zStateEstimate) ? 682:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1182 & r_state==zStateEstimate) ? 379:
			/**/
			/**/
			 /**/
			(r_counter == 1183 & r_state==zStateEstimate) ? 615:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1185 & r_state==zStateEstimate) ? 383:
			/**/
			/**/
			 /**/
			(r_counter == 1186 & r_state==zStateEstimate) ? 683:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1188 & r_state==zStateEstimate) ? 387:
			/**/
			/**/
			 /**/
			(r_counter == 1189 & r_state==zStateEstimate) ? 591:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1191 & r_state==zStateEstimate) ? 391:
			/**/
			/**/
			 /**/
			(r_counter == 1192 & r_state==zStateEstimate) ? 651:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1194 & r_state==zStateEstimate) ? 395:
			/**/
			/**/
			 /**/
			(r_counter == 1195 & r_state==zStateEstimate) ? 539:
			/**/
			/**/
			 /**/
			/**/
			 /**/
			(r_counter == 1197 & r_state==zStateEstimate) ? 399:
			/**/
			/**/
			 /**/
			(r_counter == 1198 & r_state==zStateEstimate) ? 455:
			/**/
			/**/
			 /**/
			/**/
			0;
   assign i_wdata_alpha=o_data_test_alpha;
   
   
   //beta
   assign i_wen_beta=(r_state==zStateBetaInit) | ((r_state==zStateColumn) & (
									     /**/
									     (r_counter==3) |
									     /**/
									     (r_counter==5) |
									     /**/
									     (r_counter==7) |
									     /**/
									     (r_counter==9) |
									     /**/
									     (r_counter==11) |
									     /**/
									     (r_counter==13) |
									     /**/
									     (r_counter==15) |
									     /**/
									     (r_counter==17) |
									     /**/
									     (r_counter==19) |
									     /**/
									     (r_counter==21) |
									     /**/
									     (r_counter==23) |
									     /**/
									     (r_counter==25) |
									     /**/
									     (r_counter==27) |
									     /**/
									     (r_counter==29) |
									     /**/
									     (r_counter==31) |
									     /**/
									     (r_counter==33) |
									     /**/
									     (r_counter==35) |
									     /**/
									     (r_counter==37) |
									     /**/
									     (r_counter==39) |
									     /**/
									     (r_counter==41) |
									     /**/
									     (r_counter==43) |
									     /**/
									     (r_counter==45) |
									     /**/
									     (r_counter==47) |
									     /**/
									     (r_counter==49) |
									     /**/
									     (r_counter==51) |
									     /**/
									     (r_counter==53) |
									     /**/
									     (r_counter==55) |
									     /**/
									     (r_counter==57) |
									     /**/
									     (r_counter==59) |
									     /**/
									     (r_counter==61) |
									     /**/
									     (r_counter==63) |
									     /**/
									     (r_counter==65) |
									     /**/
									     (r_counter==67) |
									     /**/
									     (r_counter==69) |
									     /**/
									     (r_counter==71) |
									     /**/
									     (r_counter==73) |
									     /**/
									     (r_counter==75) |
									     /**/
									     (r_counter==77) |
									     /**/
									     (r_counter==79) |
									     /**/
									     (r_counter==81) |
									     /**/
									     (r_counter==83) |
									     /**/
									     (r_counter==85) |
									     /**/
									     (r_counter==87) |
									     /**/
									     (r_counter==89) |
									     /**/
									     (r_counter==91) |
									     /**/
									     (r_counter==93) |
									     /**/
									     (r_counter==95) |
									     /**/
									     (r_counter==97) |
									     /**/
									     (r_counter==99) |
									     /**/
									     (r_counter==101) |
									     /**/
									     (r_counter==103) |
									     /**/
									     (r_counter==105) |
									     /**/
									     (r_counter==107) |
									     /**/
									     (r_counter==109) |
									     /**/
									     (r_counter==111) |
									     /**/
									     (r_counter==113) |
									     /**/
									     (r_counter==115) |
									     /**/
									     (r_counter==117) |
									     /**/
									     (r_counter==119) |
									     /**/
									     (r_counter==121) |
									     /**/
									     (r_counter==123) |
									     /**/
									     (r_counter==125) |
									     /**/
									     (r_counter==127) |
									     /**/
									     (r_counter==129) |
									     /**/
									     (r_counter==131) |
									     /**/
									     (r_counter==133) |
									     /**/
									     (r_counter==135) |
									     /**/
									     (r_counter==137) |
									     /**/
									     (r_counter==139) |
									     /**/
									     (r_counter==141) |
									     /**/
									     (r_counter==143) |
									     /**/
									     (r_counter==145) |
									     /**/
									     (r_counter==147) |
									     /**/
									     (r_counter==149) |
									     /**/
									     (r_counter==151) |
									     /**/
									     (r_counter==153) |
									     /**/
									     (r_counter==155) |
									     /**/
									     (r_counter==157) |
									     /**/
									     (r_counter==159) |
									     /**/
									     (r_counter==161) |
									     /**/
									     (r_counter==163) |
									     /**/
									     (r_counter==165) |
									     /**/
									     (r_counter==167) |
									     /**/
									     (r_counter==169) |
									     /**/
									     (r_counter==171) |
									     /**/
									     (r_counter==173) |
									     /**/
									     (r_counter==175) |
									     /**/
									     (r_counter==177) |
									     /**/
									     (r_counter==179) |
									     /**/
									     (r_counter==181) |
									     /**/
									     (r_counter==183) |
									     /**/
									     (r_counter==185) |
									     /**/
									     (r_counter==187) |
									     /**/
									     (r_counter==189) |
									     /**/
									     (r_counter==191) |
									     /**/
									     (r_counter==193) |
									     /**/
									     (r_counter==195) |
									     /**/
									     (r_counter==197) |
									     /**/
									     (r_counter==199) |
									     /**/
									     (r_counter==201) |
									     /**/
									     (r_counter==203) |
									     /**/
									     (r_counter==205) |
									     /**/
									     (r_counter==207) |
									     /**/
									     (r_counter==209) |
									     /**/
									     (r_counter==211) |
									     /**/
									     (r_counter==213) |
									     /**/
									     (r_counter==215) |
									     /**/
									     (r_counter==217) |
									     /**/
									     (r_counter==219) |
									     /**/
									     (r_counter==221) |
									     /**/
									     (r_counter==223) |
									     /**/
									     (r_counter==225) |
									     /**/
									     (r_counter==227) |
									     /**/
									     (r_counter==229) |
									     /**/
									     (r_counter==231) |
									     /**/
									     (r_counter==233) |
									     /**/
									     (r_counter==235) |
									     /**/
									     (r_counter==237) |
									     /**/
									     (r_counter==239) |
									     /**/
									     (r_counter==241) |
									     /**/
									     (r_counter==243) |
									     /**/
									     (r_counter==245) |
									     /**/
									     (r_counter==247) |
									     /**/
									     (r_counter==249) |
									     /**/
									     (r_counter==251) |
									     /**/
									     (r_counter==253) |
									     /**/
									     (r_counter==255) |
									     /**/
									     (r_counter==257) |
									     /**/
									     (r_counter==259) |
									     /**/
									     (r_counter==261) |
									     /**/
									     (r_counter==263) |
									     /**/
									     (r_counter==265) |
									     /**/
									     (r_counter==267) |
									     /**/
									     (r_counter==269) |
									     /**/
									     (r_counter==271) |
									     /**/
									     (r_counter==273) |
									     /**/
									     (r_counter==275) |
									     /**/
									     (r_counter==277) |
									     /**/
									     (r_counter==279) |
									     /**/
									     (r_counter==281) |
									     /**/
									     (r_counter==283) |
									     /**/
									     (r_counter==285) |
									     /**/
									     (r_counter==287) |
									     /**/
									     (r_counter==289) |
									     /**/
									     (r_counter==291) |
									     /**/
									     (r_counter==293) |
									     /**/
									     (r_counter==295) |
									     /**/
									     (r_counter==297) |
									     /**/
									     (r_counter==299) |
									     /**/
									     (r_counter==301) |
									     /**/
									     (r_counter==303) |
									     /**/
									     (r_counter==305) |
									     /**/
									     (r_counter==307) |
									     /**/
									     (r_counter==309) |
									     /**/
									     (r_counter==311) |
									     /**/
									     (r_counter==313) |
									     /**/
									     (r_counter==315) |
									     /**/
									     (r_counter==317) |
									     /**/
									     (r_counter==319) |
									     /**/
									     (r_counter==321) |
									     /**/
									     (r_counter==323) |
									     /**/
									     (r_counter==325) |
									     /**/
									     (r_counter==327) |
									     /**/
									     (r_counter==329) |
									     /**/
									     (r_counter==331) |
									     /**/
									     (r_counter==333) |
									     /**/
									     (r_counter==335) |
									     /**/
									     (r_counter==337) |
									     /**/
									     (r_counter==339) |
									     /**/
									     (r_counter==341) |
									     /**/
									     (r_counter==343) |
									     /**/
									     (r_counter==345) |
									     /**/
									     (r_counter==347) |
									     /**/
									     (r_counter==349) |
									     /**/
									     (r_counter==351) |
									     /**/
									     (r_counter==353) |
									     /**/
									     (r_counter==355) |
									     /**/
									     (r_counter==357) |
									     /**/
									     (r_counter==359) |
									     /**/
									     (r_counter==361) |
									     /**/
									     (r_counter==363) |
									     /**/
									     (r_counter==365) |
									     /**/
									     (r_counter==367) |
									     /**/
									     (r_counter==369) |
									     /**/
									     (r_counter==371) |
									     /**/
									     (r_counter==373) |
									     /**/
									     (r_counter==375) |
									     /**/
									     (r_counter==377) |
									     /**/
									     (r_counter==379) |
									     /**/
									     (r_counter==381) |
									     /**/
									     (r_counter==383) |
									     /**/
									     (r_counter==385) |
									     /**/
									     (r_counter==387) |
									     /**/
									     (r_counter==389) |
									     /**/
									     (r_counter==391) |
									     /**/
									     (r_counter==393) |
									     /**/
									     (r_counter==395) |
									     /**/
									     (r_counter==397) |
									     /**/
									     (r_counter==399) |
									     /**/
									     (r_counter==401) |
									     /**/
									     (r_counter==403) |
									     /**/
									     (r_counter==405) |
									     /**/
									     (r_counter==407) |
									     /**/
									     (r_counter==409) |
									     /**/
									     (r_counter==411) |
									     /**/
									     (r_counter==413) |
									     /**/
									     (r_counter==415) |
									     /**/
									     (r_counter==417) |
									     /**/
									     (r_counter==419) |
									     /**/
									     (r_counter==421) |
									     /**/
									     (r_counter==423) |
									     /**/
									     (r_counter==425) |
									     /**/
									     (r_counter==427) |
									     /**/
									     (r_counter==429) |
									     /**/
									     (r_counter==431) |
									     /**/
									     (r_counter==433) |
									     /**/
									     (r_counter==435) |
									     /**/
									     (r_counter==437) |
									     /**/
									     (r_counter==439) |
									     /**/
									     (r_counter==441) |
									     /**/
									     (r_counter==443) |
									     /**/
									     (r_counter==445) |
									     /**/
									     (r_counter==447) |
									     /**/
									     (r_counter==449) |
									     /**/
									     (r_counter==451) |
									     /**/
									     (r_counter==453) |
									     /**/
									     (r_counter==455) |
									     /**/
									     (r_counter==457) |
									     /**/
									     (r_counter==459) |
									     /**/
									     (r_counter==461) |
									     /**/
									     (r_counter==463) |
									     /**/
									     (r_counter==465) |
									     /**/
									     (r_counter==467) |
									     /**/
									     (r_counter==469) |
									     /**/
									     (r_counter==471) |
									     /**/
									     (r_counter==473) |
									     /**/
									     (r_counter==475) |
									     /**/
									     (r_counter==477) |
									     /**/
									     (r_counter==479) |
									     /**/
									     (r_counter==481) |
									     /**/
									     (r_counter==483) |
									     /**/
									     (r_counter==485) |
									     /**/
									     (r_counter==487) |
									     /**/
									     (r_counter==489) |
									     /**/
									     (r_counter==491) |
									     /**/
									     (r_counter==493) |
									     /**/
									     (r_counter==495) |
									     /**/
									     (r_counter==497) |
									     /**/
									     (r_counter==499) |
									     /**/
									     (r_counter==501) |
									     /**/
									     (r_counter==503) |
									     /**/
									     (r_counter==505) |
									     /**/
									     (r_counter==507) |
									     /**/
									     (r_counter==509) |
									     /**/
									     (r_counter==511) |
									     /**/
									     (r_counter==513) |
									     /**/
									     (r_counter==515) |
									     /**/
									     (r_counter==517) |
									     /**/
									     (r_counter==519) |
									     /**/
									     (r_counter==521) |
									     /**/
									     (r_counter==523) |
									     /**/
									     (r_counter==525) |
									     /**/
									     (r_counter==527) |
									     /**/
									     (r_counter==529) |
									     /**/
									     (r_counter==531) |
									     /**/
									     (r_counter==533) |
									     /**/
									     (r_counter==535) |
									     /**/
									     (r_counter==537) |
									     /**/
									     (r_counter==539) |
									     /**/
									     (r_counter==541) |
									     /**/
									     (r_counter==543) |
									     /**/
									     (r_counter==545) |
									     /**/
									     (r_counter==547) |
									     /**/
									     (r_counter==549) |
									     /**/
									     (r_counter==551) |
									     /**/
									     (r_counter==553) |
									     /**/
									     (r_counter==555) |
									     /**/
									     (r_counter==557) |
									     /**/
									     (r_counter==559) |
									     /**/
									     (r_counter==561) |
									     /**/
									     (r_counter==563) |
									     /**/
									     (r_counter==565) |
									     /**/
									     (r_counter==567) |
									     /**/
									     (r_counter==569) |
									     /**/
									     (r_counter==571) |
									     /**/
									     (r_counter==573) |
									     /**/
									     (r_counter==575) |
									     /**/
									     (r_counter==577) |
									     /**/
									     (r_counter==579) |
									     /**/
									     (r_counter==581) |
									     /**/
									     (r_counter==583) |
									     /**/
									     (r_counter==585) |
									     /**/
									     (r_counter==587) |
									     /**/
									     (r_counter==589) |
									     /**/
									     (r_counter==591) |
									     /**/
									     (r_counter==593) |
									     /**/
									     (r_counter==595) |
									     /**/
									     (r_counter==597) |
									     /**/
									     (r_counter==599) |
									     /**/
									     (r_counter==601) |
									     /**/
									     (r_counter==603) |
									     /**/
									     (r_counter==605) |
									     /**/
									     (r_counter==607) |
									     /**/
									     (r_counter==609) |
									     /**/
									     (r_counter==611) |
									     /**/
									     (r_counter==613) |
									     /**/
									     (r_counter==615) |
									     /**/
									     (r_counter==617) |
									     /**/
									     (r_counter==619) |
									     /**/
									     (r_counter==621) |
									     /**/
									     (r_counter==623) |
									     /**/
									     (r_counter==625) |
									     /**/
									     (r_counter==627) |
									     /**/
									     (r_counter==629) |
									     /**/
									     (r_counter==631) |
									     /**/
									     (r_counter==633) |
									     /**/
									     (r_counter==635) |
									     /**/
									     (r_counter==637) |
									     /**/
									     (r_counter==639) |
									     /**/
									     (r_counter==641) |
									     /**/
									     (r_counter==643) |
									     /**/
									     (r_counter==645) |
									     /**/
									     (r_counter==647) |
									     /**/
									     (r_counter==649) |
									     /**/
									     (r_counter==651) |
									     /**/
									     (r_counter==653) |
									     /**/
									     (r_counter==655) |
									     /**/
									     (r_counter==657) |
									     /**/
									     (r_counter==659) |
									     /**/
									     (r_counter==661) |
									     /**/
									     (r_counter==663) |
									     /**/
									     (r_counter==665) |
									     /**/
									     (r_counter==667) |
									     /**/
									     (r_counter==669) |
									     /**/
									     (r_counter==671) |
									     /**/
									     (r_counter==673) |
									     /**/
									     (r_counter==675) |
									     /**/
									     (r_counter==677) |
									     /**/
									     (r_counter==679) |
									     /**/
									     (r_counter==681) |
									     /**/
									     (r_counter==683) |
									     /**/
									     (r_counter==685) |
									     /**/
									     (r_counter==687) |
									     /**/
									     (r_counter==689) |
									     /**/
									     (r_counter==691) |
									     /**/
									     (r_counter==693) |
									     /**/
									     (r_counter==695) |
									     /**/
									     (r_counter==697) |
									     /**/
									     (r_counter==699) |
									     /**/
									     (r_counter==701) |
									     /**/
									     (r_counter==703) |
									     /**/
									     (r_counter==705) |
									     /**/
									     (r_counter==707) |
									     /**/
									     (r_counter==709) |
									     /**/
									     (r_counter==711) |
									     /**/
									     (r_counter==713) |
									     /**/
									     (r_counter==715) |
									     /**/
									     (r_counter==717) |
									     /**/
									     (r_counter==719) |
									     /**/
									     (r_counter==721) |
									     /**/
									     (r_counter==723) |
									     /**/
									     (r_counter==725) |
									     /**/
									     (r_counter==727) |
									     /**/
									     (r_counter==729) |
									     /**/
									     (r_counter==731) |
									     /**/
									     (r_counter==733) |
									     /**/
									     (r_counter==735) |
									     /**/
									     (r_counter==737) |
									     /**/
									     (r_counter==739) |
									     /**/
									     (r_counter==741) |
									     /**/
									     (r_counter==743) |
									     /**/
									     (r_counter==745) |
									     /**/
									     (r_counter==747) |
									     /**/
									     (r_counter==749) |
									     /**/
									     (r_counter==751) |
									     /**/
									     (r_counter==753) |
									     /**/
									     (r_counter==755) |
									     /**/
									     (r_counter==757) |
									     /**/
									     (r_counter==759) |
									     /**/
									     (r_counter==761) |
									     /**/
									     (r_counter==763) |
									     /**/
									     (r_counter==765) |
									     /**/
									     (r_counter==767) |
									     /**/
									     (r_counter==769) |
									     /**/
									     (r_counter==771) |
									     /**/
									     (r_counter==773) |
									     /**/
									     (r_counter==775) |
									     /**/
									     (r_counter==777) |
									     /**/
									     (r_counter==779) |
									     /**/
									     (r_counter==781) |
									     /**/
									     (r_counter==783) |
									     /**/
									     (r_counter==785) |
									     /**/
									     (r_counter==787) |
									     /**/
									     (r_counter==789) |
									     /**/
									     (r_counter==791) |
									     /**/
									     (r_counter==793) |
									     /**/
									     (r_counter==795) |
									     /**/
									     (r_counter==797) |
									     /**/
									     (r_counter==799) |
									     /**/
									     (r_counter==801) |
									     /**/
									     (r_counter==803) |
									     /**/
									     (r_counter==805) |
									     /**/
									     (r_counter==807) |
									     /**/
									     (r_counter==809) |
									     /**/
									     (r_counter==811) |
									     /**/
									     (r_counter==813) |
									     /**/
									     (r_counter==815) |
									     /**/
									     (r_counter==817) |
									     /**/
									     (r_counter==819) |
									     /**/
									     (r_counter==821) |
									     /**/
									     (r_counter==823) |
									     /**/
									     (r_counter==825) |
									     /**/
									     (r_counter==827) |
									     /**/
									     (r_counter==829) |
									     /**/
									     (r_counter==831) |
									     /**/
									     (r_counter==833) |
									     /**/
									     (r_counter==835) |
									     /**/
									     (r_counter==837) |
									     /**/
									     (r_counter==839) |
									     /**/
									     (r_counter==841) |
									     /**/
									     (r_counter==843) |
									     /**/
									     (r_counter==845) |
									     /**/
									     (r_counter==847) |
									     /**/
									     (r_counter==849) |
									     /**/
									     (r_counter==851) |
									     /**/
									     (r_counter==853) |
									     /**/
									     (r_counter==855) |
									     /**/
									     (r_counter==857) |
									     /**/
									     (r_counter==859) |
									     /**/
									     (r_counter==861) |
									     /**/
									     (r_counter==863) |
									     /**/
									     (r_counter==865) |
									     /**/
									     (r_counter==867) |
									     /**/
									     (r_counter==869) |
									     /**/
									     (r_counter==871) |
									     /**/
									     (r_counter==873) |
									     /**/
									     (r_counter==875) |
									     /**/
									     (r_counter==877) |
									     /**/
									     (r_counter==879) |
									     /**/
									     (r_counter==881) |
									     /**/
									     (r_counter==883) |
									     /**/
									     (r_counter==885) |
									     /**/
									     (r_counter==887) |
									     /**/
									     (r_counter==889) |
									     /**/
									     (r_counter==891) |
									     /**/
									     (r_counter==893) |
									     /**/
									     (r_counter==895) |
									     /**/
									     (r_counter==897) |
									     /**/
									     (r_counter==899) |
									     /**/
									     (r_counter==901) |
									     /**/
									     (r_counter==903) |
									     /**/
									     (r_counter==905) |
									     /**/
									     (r_counter==907) |
									     /**/
									     (r_counter==909) |
									     /**/
									     (r_counter==911) |
									     /**/
									     (r_counter==913) |
									     /**/
									     (r_counter==915) |
									     /**/
									     (r_counter==917) |
									     /**/
									     (r_counter==919) |
									     /**/
									     (r_counter==921) |
									     /**/
									     (r_counter==923) |
									     /**/
									     (r_counter==925) |
									     /**/
									     (r_counter==927) |
									     /**/
									     (r_counter==929) |
									     /**/
									     (r_counter==931) |
									     /**/
									     (r_counter==933) |
									     /**/
									     (r_counter==935) |
									     /**/
									     (r_counter==937) |
									     /**/
									     (r_counter==939) |
									     /**/
									     (r_counter==941) |
									     /**/
									     (r_counter==943) |
									     /**/
									     (r_counter==945) |
									     /**/
									     (r_counter==947) |
									     /**/
									     (r_counter==949) |
									     /**/
									     (r_counter==951) |
									     /**/
									     (r_counter==953) |
									     /**/
									     (r_counter==955) |
									     /**/
									     (r_counter==957) |
									     /**/
									     (r_counter==959) |
									     /**/
									     (r_counter==961) |
									     /**/
									     (r_counter==963) |
									     /**/
									     (r_counter==965) |
									     /**/
									     (r_counter==967) |
									     /**/
									     (r_counter==969) |
									     /**/
									     (r_counter==971) |
									     /**/
									     (r_counter==973) |
									     /**/
									     (r_counter==975) |
									     /**/
									     (r_counter==977) |
									     /**/
									     (r_counter==979) |
									     /**/
									     (r_counter==981) |
									     /**/
									     (r_counter==983) |
									     /**/
									     (r_counter==985) |
									     /**/
									     (r_counter==987) |
									     /**/
									     (r_counter==989) |
									     /**/
									     (r_counter==991) |
									     /**/
									     (r_counter==993) |
									     /**/
									     (r_counter==995) |
									     /**/
									     (r_counter==997) |
									     /**/
									     (r_counter==999) |
									     /**/
									     (r_counter==1001) |
									     /**/
									     (r_counter==1003) |
									     /**/
									     (r_counter==1005) |
									     /**/
									     (r_counter==1007) |
									     /**/
									     (r_counter==1009) |
									     /**/
									     (r_counter==1011) |
									     /**/
									     (r_counter==1013) |
									     /**/
									     (r_counter==1015) |
									     /**/
									     (r_counter==1017) |
									     /**/
									     (r_counter==1019) |
									     /**/
									     (r_counter==1021) |
									     /**/
									     (r_counter==1023) |
									     /**/
									     (r_counter==1025) |
									     /**/
									     (r_counter==1027) |
									     /**/
									     (r_counter==1029) |
									     /**/
									     (r_counter==1031) |
									     /**/
									     (r_counter==1033) |
									     /**/
									     (r_counter==1035) |
									     /**/
									     (r_counter==1037) |
									     /**/
									     (r_counter==1039) |
									     /**/
									     (r_counter==1041) |
									     /**/
									     (r_counter==1043) |
									     /**/
									     (r_counter==1045) |
									     /**/
									     (r_counter==1047) |
									     /**/
									     (r_counter==1049) |
									     /**/
									     (r_counter==1051) |
									     /**/
									     (r_counter==1053) |
									     /**/
									     (r_counter==1055) |
									     /**/
									     (r_counter==1057) |
									     /**/
									     (r_counter==1059) |
									     /**/
									     (r_counter==1061) |
									     /**/
									     (r_counter==1063) |
									     /**/
									     (r_counter==1065) |
									     /**/
									     (r_counter==1067) |
									     /**/
									     (r_counter==1069) |
									     /**/
									     (r_counter==1071) |
									     /**/
									     (r_counter==1073) |
									     /**/
									     (r_counter==1075) |
									     /**/
									     (r_counter==1077) |
									     /**/
									     (r_counter==1079) |
									     /**/
									     (r_counter==1081) |
									     /**/
									     (r_counter==1083) |
									     /**/
									     (r_counter==1085) |
									     /**/
									     (r_counter==1087) |
									     /**/
									     (r_counter==1089) |
									     /**/
									     (r_counter==1091) |
									     /**/
									     (r_counter==1093) |
									     /**/
									     (r_counter==1095) |
									     /**/
									     (r_counter==1097) |
									     /**/
									     (r_counter==1099) |
									     /**/
									     (r_counter==1101) |
									     /**/
									     (r_counter==1103) |
									     /**/
									     (r_counter==1105) |
									     /**/
									     (r_counter==1107) |
									     /**/
									     (r_counter==1109) |
									     /**/
									     (r_counter==1111) |
									     /**/
									     (r_counter==1113) |
									     /**/
									     (r_counter==1115) |
									     /**/
									     (r_counter==1117) |
									     /**/
									     (r_counter==1119) |
									     /**/
									     (r_counter==1121) |
									     /**/
									     (r_counter==1123) |
									     /**/
									     (r_counter==1125) |
									     /**/
									     (r_counter==1127) |
									     /**/
									     (r_counter==1129) |
									     /**/
									     (r_counter==1131) |
									     /**/
									     (r_counter==1133) |
									     /**/
									     (r_counter==1135) |
									     /**/
									     (r_counter==1137) |
									     /**/
									     (r_counter==1139) |
									     /**/
									     (r_counter==1141) |
									     /**/
									     (r_counter==1143) |
									     /**/
									     (r_counter==1145) |
									     /**/
									     (r_counter==1147) |
									     /**/
									     (r_counter==1149) |
									     /**/
									     (r_counter==1151) |
									     /**/
									     (r_counter==1153) |
									     /**/
									     (r_counter==1155) |
									     /**/
									     (r_counter==1157) |
									     /**/
									     (r_counter==1159) |
									     /**/
									     (r_counter==1161) |
									     /**/
									     (r_counter==1163) |
									     /**/
									     (r_counter==1165) |
									     /**/
									     (r_counter==1167) |
									     /**/
									     (r_counter==1169) |
									     /**/
									     (r_counter==1171) |
									     /**/
									     (r_counter==1173) |
									     /**/
									     (r_counter==1175) |
									     /**/
									     (r_counter==1177) |
									     /**/
									     (r_counter==1179) |
									     /**/
									     (r_counter==1181) |
									     /**/
									     (r_counter==1183) |
									     /**/
									     (r_counter==1185) |
									     /**/
									     (r_counter==1187) |
									     /**/
									     (r_counter==1189) |
									     /**/
									     (r_counter==1191) |
									     /**/
									     (r_counter==1193) |
									     /**/
									     (r_counter==1195) |
									     /**/
									     (r_counter==1197) |
									     /**/
									     (r_counter==1199) |
									     /**/
									     (r_counter==1201) |
									     /**/
									     (r_counter==1203) |
									     /**/
									     (r_counter==1205) |
									     /**/
									     (r_counter==1207) |
									     /**/
									     (r_counter==1209) |
									     /**/
									     (r_counter==1211) |
									     /**/
									     (r_counter==1213) |
									     /**/
									     (r_counter==1215) |
									     /**/
									     (r_counter==1217) |
									     /**/
									     (r_counter==1219) |
									     /**/
									     (r_counter==1221) |
									     /**/
									     (r_counter==1223) |
									     /**/
									     (r_counter==1225) |
									     /**/
									     (r_counter==1227) |
									     /**/
									     (r_counter==1229) |
									     /**/
									     (r_counter==1231) |
									     /**/
									     (r_counter==1233) |
									     /**/
									     (r_counter==1235) |
									     /**/
									     (r_counter==1237) |
									     /**/
									     (r_counter==1239) |
									     /**/
									     (r_counter==1241) |
									     /**/
									     (r_counter==1243) |
									     /**/
									     (r_counter==1245) |
									     /**/
									     (r_counter==1247) |
									     /**/
									     (r_counter==1249) |
									     /**/
									     (r_counter==1251) |
									     /**/
									     (r_counter==1253) |
									     /**/
									     (r_counter==1255) |
									     /**/
									     (r_counter==1257) |
									     /**/
									     (r_counter==1259) |
									     /**/
									     (r_counter==1261) |
									     /**/
									     (r_counter==1263) |
									     /**/
									     (r_counter==1265) |
									     /**/
									     (r_counter==1267) |
									     /**/
									     (r_counter==1269) |
									     /**/
									     (r_counter==1271) |
									     /**/
									     (r_counter==1273) |
									     /**/
									     (r_counter==1275) |
									     /**/
									     (r_counter==1277) |
									     /**/
									     (r_counter==1279) |
									     /**/
									     (r_counter==1281) |
									     /**/
									     (r_counter==1283) |
									     /**/
									     (r_counter==1285) |
									     /**/
									     (r_counter==1287) |
									     /**/
									     (r_counter==1289) |
									     /**/
									     (r_counter==1291) |
									     /**/
									     (r_counter==1293) |
									     /**/
									     (r_counter==1295) |
									     /**/
									     (r_counter==1297) |
									     /**/
									     (r_counter==1299) |
									     /**/
									     (r_counter==1301) |
									     /**/
									     (r_counter==1303) |
									     /**/
									     (r_counter==1305) |
									     /**/
									     (r_counter==1307) |
									     /**/
									     (r_counter==1309) |
									     /**/
									     (r_counter==1311) |
									     /**/
									     (r_counter==1313) |
									     /**/
									     (r_counter==1315) |
									     /**/
									     (r_counter==1317) |
									     /**/
									     (r_counter==1319) |
									     /**/
									     (r_counter==1321) |
									     /**/
									     (r_counter==1323) |
									     /**/
									     (r_counter==1325) |
									     /**/
									     (r_counter==1327) |
									     /**/
									     (r_counter==1329) |
									     /**/
									     (r_counter==1331) |
									     /**/
									     (r_counter==1333) |
									     /**/
									     (r_counter==1335) |
									     /**/
									     (r_counter==1337) |
									     /**/
									     (r_counter==1339) |
									     /**/
									     (r_counter==1341) |
									     /**/
									     (r_counter==1343) |
									     /**/
									     (r_counter==1345) |
									     /**/
									     (r_counter==1347) |
									     /**/
									     (r_counter==1349) |
									     /**/
									     (r_counter==1351) |
									     /**/
									     (r_counter==1353) |
									     /**/
									     (r_counter==1355) |
									     /**/
									     (r_counter==1357) |
									     /**/
									     (r_counter==1359) |
									     /**/
									     (r_counter==1361) |
									     /**/
									     (r_counter==1363) |
									     /**/
									     (r_counter==1365) |
									     /**/
									     (r_counter==1367) |
									     /**/
									     (r_counter==1369) |
									     /**/
									     (r_counter==1371) |
									     /**/
									     (r_counter==1373) |
									     /**/
									     (r_counter==1375) |
									     /**/
									     (r_counter==1377) |
									     /**/
									     (r_counter==1379) |
									     /**/
									     (r_counter==1381) |
									     /**/
									     (r_counter==1383) |
									     /**/
									     (r_counter==1385) |
									     /**/
									     (r_counter==1387) |
									     /**/
									     (r_counter==1389) |
									     /**/
									     (r_counter==1391) |
									     /**/
									     (r_counter==1393) |
									     /**/
									     (r_counter==1395) |
									     /**/
									     (r_counter==1397) |
									     /**/
									     (r_counter==1399) |
									     /**/
									     (r_counter==1401) |
									     /**/
									     (r_counter==1403) |
									     /**/
									     (r_counter==1405) |
									     /**/
									     (r_counter==1407) |
									     /**/
									     (r_counter==1409) |
									     /**/
									     (r_counter==1411) |
									     /**/
									     (r_counter==1413) |
									     /**/
									     (r_counter==1415) |
									     /**/
									     (r_counter==1417) |
									     /**/
									     (r_counter==1419) |
									     /**/
									     (r_counter==1421) |
									     /**/
									     (r_counter==1423) |
									     /**/
									     (r_counter==1425) |
									     /**/
									     (r_counter==1427) |
									     /**/
									     (r_counter==1429) |
									     /**/
									     (r_counter==1431) |
									     /**/
									     (r_counter==1433) |
									     /**/
									     (r_counter==1435) |
									     /**/
									     (r_counter==1437) |
									     /**/
									     (r_counter==1439) |
									     /**/
									     (r_counter==1441) |
									     /**/
									     (r_counter==1443) |
									     /**/
									     (r_counter==1445) |
									     /**/
									     (r_counter==1447) |
									     /**/
									     (r_counter==1449) |
									     /**/
									     (r_counter==1451) |
									     /**/
									     (r_counter==1453) |
									     /**/
									     (r_counter==1455) |
									     /**/
									     (r_counter==1457) |
									     /**/
									     (r_counter==1459) |
									     /**/
									     (r_counter==1461) |
									     /**/
									     (r_counter==1463) |
									     /**/
									     (r_counter==1465) |
									     /**/
									     (r_counter==1467) |
									     /**/
									     (r_counter==1469) |
									     /**/
									     (r_counter==1471) |
									     /**/
									     (r_counter==1473) |
									     /**/
									     (r_counter==1475) |
									     /**/
									     (r_counter==1477) |
									     /**/
									     (r_counter==1479) |
									     /**/
									     (r_counter==1481) |
									     /**/
									     (r_counter==1483) |
									     /**/
									     (r_counter==1485) |
									     /**/
									     (r_counter==1487) |
									     /**/
									     (r_counter==1489) |
									     /**/
									     (r_counter==1491) |
									     /**/
									     (r_counter==1493) |
									     /**/
									     (r_counter==1495) |
									     /**/
									     (r_counter==1497) |
									     /**/
									     (r_counter==1499) |
									     /**/
									     (r_counter==1501) |
									     /**/
									     (r_counter==1503) |
									     /**/
									     (r_counter==1505) |
									     /**/
									     (r_counter==1507) |
									     /**/
									     (r_counter==1509) |
									     /**/
									     (r_counter==1511) |
									     /**/
									     (r_counter==1513) |
									     /**/
									     (r_counter==1515) |
									     /**/
									     (r_counter==1517) |
									     /**/
									     (r_counter==1519) |
									     /**/
									     (r_counter==1521) |
									     /**/
									     (r_counter==1523) |
									     /**/
									     (r_counter==1525) |
									     /**/
									     (r_counter==1527) |
									     /**/
									     (r_counter==1529) |
									     /**/
									     (r_counter==1531) |
									     /**/
									     (r_counter==1533) |
									     /**/
									     (r_counter==1535) |
									     /**/
									     (r_counter==1537) |
									     /**/
									     (r_counter==1539) |
									     /**/
									     (r_counter==1541) |
									     /**/
									     (r_counter==1543) |
									     /**/
									     (r_counter==1545) |
									     /**/
									     (r_counter==1547) |
									     /**/
									     (r_counter==1549) |
									     /**/
									     (r_counter==1551) |
									     /**/
									     (r_counter==1553) |
									     /**/
									     (r_counter==1555) |
									     /**/
									     (r_counter==1557) |
									     /**/
									     (r_counter==1559) |
									     /**/
									     (r_counter==1561) |
									     /**/
									     (r_counter==1563) |
									     /**/
									     (r_counter==1565) |
									     /**/
									     (r_counter==1567) |
									     /**/
									     (r_counter==1569) |
									     /**/
									     (r_counter==1571) |
									     /**/
									     (r_counter==1573) |
									     /**/
									     (r_counter==1575) |
									     /**/
									     (r_counter==1577) |
									     /**/
									     (r_counter==1579) |
									     /**/
									     (r_counter==1581) |
									     /**/
									     (r_counter==1583) |
									     /**/
									     (r_counter==1585) |
									     /**/
									     (r_counter==1587) |
									     /**/
									     (r_counter==1589) |
									     /**/
									     (r_counter==1591) |
									     /**/
									     (r_counter==1593) |
									     /**/
									     (r_counter==1595) |
									     /**/
									     (r_counter==1597) |
									     /**/
									     (r_counter==1599) |
									     /**/
									     (r_counter==1601)));
   
   assign i_waddr_beta=(r_state == zStateBetaInit & r_counter!=0) ? r_counter-1:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 3) ? 0:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 5) ? 1:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 7) ? 2:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 9) ? 3:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 11) ? 4:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 13) ? 5:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 15) ? 6:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 17) ? 7:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 19) ? 8:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 21) ? 9:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 23) ? 10:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 25) ? 11:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 27) ? 12:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 29) ? 13:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 31) ? 14:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 33) ? 15:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 35) ? 16:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 37) ? 17:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 39) ? 18:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 41) ? 19:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 43) ? 20:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 45) ? 21:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 47) ? 22:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 49) ? 23:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 51) ? 24:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 53) ? 25:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 55) ? 26:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 57) ? 27:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 59) ? 28:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 61) ? 29:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 63) ? 30:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 65) ? 31:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 67) ? 32:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 69) ? 33:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 71) ? 34:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 73) ? 35:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 75) ? 36:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 77) ? 37:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 79) ? 38:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 81) ? 39:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 83) ? 40:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 85) ? 41:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 87) ? 42:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 89) ? 43:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 91) ? 44:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 93) ? 45:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 95) ? 46:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 97) ? 47:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 99) ? 48:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 101) ? 49:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 103) ? 50:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 105) ? 51:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 107) ? 52:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 109) ? 53:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 111) ? 54:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 113) ? 55:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 115) ? 56:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 117) ? 57:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 119) ? 58:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 121) ? 59:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 123) ? 60:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 125) ? 61:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 127) ? 62:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 129) ? 63:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 131) ? 64:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 133) ? 65:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 135) ? 66:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 137) ? 67:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 139) ? 68:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 141) ? 69:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 143) ? 70:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 145) ? 71:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 147) ? 72:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 149) ? 73:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 151) ? 74:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 153) ? 75:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 155) ? 76:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 157) ? 77:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 159) ? 78:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 161) ? 79:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 163) ? 80:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 165) ? 81:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 167) ? 82:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 169) ? 83:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 171) ? 84:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 173) ? 85:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 175) ? 86:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 177) ? 87:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 179) ? 88:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 181) ? 89:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 183) ? 90:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 185) ? 91:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 187) ? 92:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 189) ? 93:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 191) ? 94:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 193) ? 95:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 195) ? 96:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 197) ? 97:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 199) ? 98:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 201) ? 99:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 203) ? 100:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 205) ? 101:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 207) ? 102:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 209) ? 103:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 211) ? 104:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 213) ? 105:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 215) ? 106:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 217) ? 107:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 219) ? 108:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 221) ? 109:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 223) ? 110:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 225) ? 111:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 227) ? 112:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 229) ? 113:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 231) ? 114:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 233) ? 115:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 235) ? 116:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 237) ? 117:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 239) ? 118:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 241) ? 119:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 243) ? 120:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 245) ? 121:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 247) ? 122:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 249) ? 123:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 251) ? 124:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 253) ? 125:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 255) ? 126:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 257) ? 127:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 259) ? 128:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 261) ? 129:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 263) ? 130:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 265) ? 131:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 267) ? 132:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 269) ? 133:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 271) ? 134:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 273) ? 135:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 275) ? 136:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 277) ? 137:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 279) ? 138:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 281) ? 139:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 283) ? 140:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 285) ? 141:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 287) ? 142:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 289) ? 143:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 291) ? 144:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 293) ? 145:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 295) ? 146:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 297) ? 147:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 299) ? 148:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 301) ? 149:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 303) ? 150:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 305) ? 151:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 307) ? 152:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 309) ? 153:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 311) ? 154:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 313) ? 155:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 315) ? 156:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 317) ? 157:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 319) ? 158:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 321) ? 159:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 323) ? 160:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 325) ? 161:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 327) ? 162:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 329) ? 163:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 331) ? 164:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 333) ? 165:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 335) ? 166:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 337) ? 167:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 339) ? 168:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 341) ? 169:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 343) ? 170:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 345) ? 171:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 347) ? 172:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 349) ? 173:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 351) ? 174:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 353) ? 175:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 355) ? 176:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 357) ? 177:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 359) ? 178:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 361) ? 179:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 363) ? 180:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 365) ? 181:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 367) ? 182:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 369) ? 183:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 371) ? 184:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 373) ? 185:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 375) ? 186:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 377) ? 187:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 379) ? 188:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 381) ? 189:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 383) ? 190:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 385) ? 191:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 387) ? 192:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 389) ? 193:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 391) ? 194:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 393) ? 195:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 395) ? 196:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 397) ? 197:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 399) ? 198:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 401) ? 199:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 403) ? 200:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 405) ? 201:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 407) ? 202:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 409) ? 203:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 411) ? 204:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 413) ? 205:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 415) ? 206:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 417) ? 207:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 419) ? 208:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 421) ? 209:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 423) ? 210:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 425) ? 211:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 427) ? 212:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 429) ? 213:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 431) ? 214:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 433) ? 215:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 435) ? 216:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 437) ? 217:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 439) ? 218:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 441) ? 219:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 443) ? 220:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 445) ? 221:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 447) ? 222:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 449) ? 223:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 451) ? 224:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 453) ? 225:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 455) ? 226:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 457) ? 227:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 459) ? 228:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 461) ? 229:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 463) ? 230:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 465) ? 231:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 467) ? 232:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 469) ? 233:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 471) ? 234:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 473) ? 235:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 475) ? 236:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 477) ? 237:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 479) ? 238:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 481) ? 239:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 483) ? 240:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 485) ? 241:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 487) ? 242:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 489) ? 243:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 491) ? 244:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 493) ? 245:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 495) ? 246:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 497) ? 247:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 499) ? 248:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 501) ? 249:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 503) ? 250:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 505) ? 251:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 507) ? 252:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 509) ? 253:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 511) ? 254:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 513) ? 255:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 515) ? 256:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 517) ? 257:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 519) ? 258:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 521) ? 259:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 523) ? 260:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 525) ? 261:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 527) ? 262:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 529) ? 263:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 531) ? 264:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 533) ? 265:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 535) ? 266:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 537) ? 267:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 539) ? 268:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 541) ? 269:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 543) ? 270:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 545) ? 271:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 547) ? 272:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 549) ? 273:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 551) ? 274:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 553) ? 275:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 555) ? 276:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 557) ? 277:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 559) ? 278:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 561) ? 279:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 563) ? 280:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 565) ? 281:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 567) ? 282:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 569) ? 283:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 571) ? 284:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 573) ? 285:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 575) ? 286:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 577) ? 287:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 579) ? 288:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 581) ? 289:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 583) ? 290:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 585) ? 291:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 587) ? 292:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 589) ? 293:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 591) ? 294:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 593) ? 295:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 595) ? 296:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 597) ? 297:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 599) ? 298:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 601) ? 299:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 603) ? 300:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 605) ? 301:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 607) ? 302:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 609) ? 303:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 611) ? 304:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 613) ? 305:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 615) ? 306:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 617) ? 307:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 619) ? 308:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 621) ? 309:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 623) ? 310:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 625) ? 311:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 627) ? 312:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 629) ? 313:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 631) ? 314:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 633) ? 315:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 635) ? 316:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 637) ? 317:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 639) ? 318:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 641) ? 319:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 643) ? 320:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 645) ? 321:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 647) ? 322:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 649) ? 323:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 651) ? 324:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 653) ? 325:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 655) ? 326:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 657) ? 327:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 659) ? 328:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 661) ? 329:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 663) ? 330:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 665) ? 331:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 667) ? 332:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 669) ? 333:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 671) ? 334:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 673) ? 335:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 675) ? 336:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 677) ? 337:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 679) ? 338:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 681) ? 339:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 683) ? 340:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 685) ? 341:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 687) ? 342:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 689) ? 343:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 691) ? 344:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 693) ? 345:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 695) ? 346:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 697) ? 347:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 699) ? 348:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 701) ? 349:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 703) ? 350:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 705) ? 351:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 707) ? 352:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 709) ? 353:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 711) ? 354:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 713) ? 355:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 715) ? 356:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 717) ? 357:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 719) ? 358:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 721) ? 359:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 723) ? 360:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 725) ? 361:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 727) ? 362:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 729) ? 363:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 731) ? 364:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 733) ? 365:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 735) ? 366:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 737) ? 367:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 739) ? 368:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 741) ? 369:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 743) ? 370:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 745) ? 371:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 747) ? 372:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 749) ? 373:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 751) ? 374:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 753) ? 375:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 755) ? 376:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 757) ? 377:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 759) ? 378:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 761) ? 379:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 763) ? 380:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 765) ? 381:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 767) ? 382:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 769) ? 383:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 771) ? 384:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 773) ? 385:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 775) ? 386:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 777) ? 387:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 779) ? 388:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 781) ? 389:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 783) ? 390:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 785) ? 391:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 787) ? 392:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 789) ? 393:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 791) ? 394:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 793) ? 395:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 795) ? 396:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 797) ? 397:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 799) ? 398:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 801) ? 399:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 803) ? 400:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 805) ? 401:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 807) ? 402:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 809) ? 403:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 811) ? 404:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 813) ? 405:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 815) ? 406:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 817) ? 407:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 819) ? 408:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 821) ? 409:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 823) ? 410:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 825) ? 411:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 827) ? 412:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 829) ? 413:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 831) ? 414:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 833) ? 415:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 835) ? 416:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 837) ? 417:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 839) ? 418:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 841) ? 419:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 843) ? 420:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 845) ? 421:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 847) ? 422:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 849) ? 423:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 851) ? 424:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 853) ? 425:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 855) ? 426:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 857) ? 427:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 859) ? 428:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 861) ? 429:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 863) ? 430:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 865) ? 431:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 867) ? 432:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 869) ? 433:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 871) ? 434:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 873) ? 435:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 875) ? 436:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 877) ? 437:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 879) ? 438:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 881) ? 439:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 883) ? 440:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 885) ? 441:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 887) ? 442:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 889) ? 443:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 891) ? 444:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 893) ? 445:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 895) ? 446:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 897) ? 447:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 899) ? 448:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 901) ? 449:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 903) ? 450:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 905) ? 451:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 907) ? 452:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 909) ? 453:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 911) ? 454:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 913) ? 455:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 915) ? 456:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 917) ? 457:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 919) ? 458:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 921) ? 459:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 923) ? 460:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 925) ? 461:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 927) ? 462:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 929) ? 463:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 931) ? 464:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 933) ? 465:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 935) ? 466:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 937) ? 467:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 939) ? 468:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 941) ? 469:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 943) ? 470:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 945) ? 471:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 947) ? 472:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 949) ? 473:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 951) ? 474:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 953) ? 475:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 955) ? 476:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 957) ? 477:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 959) ? 478:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 961) ? 479:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 963) ? 480:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 965) ? 481:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 967) ? 482:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 969) ? 483:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 971) ? 484:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 973) ? 485:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 975) ? 486:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 977) ? 487:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 979) ? 488:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 981) ? 489:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 983) ? 490:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 985) ? 491:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 987) ? 492:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 989) ? 493:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 991) ? 494:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 993) ? 495:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 995) ? 496:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 997) ? 497:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 999) ? 498:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1001) ? 499:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1003) ? 500:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1005) ? 501:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1007) ? 502:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1009) ? 503:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1011) ? 504:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1013) ? 505:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1015) ? 506:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1017) ? 507:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1019) ? 508:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1021) ? 509:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1023) ? 510:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1025) ? 511:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1027) ? 512:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1029) ? 513:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1031) ? 514:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1033) ? 515:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1035) ? 516:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1037) ? 517:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1039) ? 518:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1041) ? 519:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1043) ? 520:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1045) ? 521:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1047) ? 522:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1049) ? 523:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1051) ? 524:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1053) ? 525:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1055) ? 526:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1057) ? 527:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1059) ? 528:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1061) ? 529:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1063) ? 530:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1065) ? 531:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1067) ? 532:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1069) ? 533:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1071) ? 534:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1073) ? 535:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1075) ? 536:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1077) ? 537:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1079) ? 538:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1081) ? 539:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1083) ? 540:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1085) ? 541:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1087) ? 542:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1089) ? 543:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1091) ? 544:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1093) ? 545:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1095) ? 546:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1097) ? 547:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1099) ? 548:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1101) ? 549:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1103) ? 550:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1105) ? 551:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1107) ? 552:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1109) ? 553:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1111) ? 554:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1113) ? 555:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1115) ? 556:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1117) ? 557:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1119) ? 558:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1121) ? 559:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1123) ? 560:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1125) ? 561:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1127) ? 562:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1129) ? 563:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1131) ? 564:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1133) ? 565:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1135) ? 566:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1137) ? 567:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1139) ? 568:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1141) ? 569:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1143) ? 570:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1145) ? 571:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1147) ? 572:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1149) ? 573:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1151) ? 574:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1153) ? 575:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1155) ? 576:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1157) ? 577:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1159) ? 578:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1161) ? 579:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1163) ? 580:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1165) ? 581:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1167) ? 582:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1169) ? 583:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1171) ? 584:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1173) ? 585:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1175) ? 586:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1177) ? 587:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1179) ? 588:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1181) ? 589:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1183) ? 590:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1185) ? 591:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1187) ? 592:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1189) ? 593:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1191) ? 594:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1193) ? 595:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1195) ? 596:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1197) ? 597:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1199) ? 598:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1201) ? 599:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1203) ? 600:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1205) ? 601:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1207) ? 602:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1209) ? 603:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1211) ? 604:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1213) ? 605:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1215) ? 606:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1217) ? 607:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1219) ? 608:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1221) ? 609:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1223) ? 610:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1225) ? 611:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1227) ? 612:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1229) ? 613:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1231) ? 614:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1233) ? 615:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1235) ? 616:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1237) ? 617:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1239) ? 618:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1241) ? 619:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1243) ? 620:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1245) ? 621:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1247) ? 622:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1249) ? 623:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1251) ? 624:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1253) ? 625:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1255) ? 626:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1257) ? 627:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1259) ? 628:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1261) ? 629:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1263) ? 630:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1265) ? 631:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1267) ? 632:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1269) ? 633:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1271) ? 634:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1273) ? 635:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1275) ? 636:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1277) ? 637:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1279) ? 638:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1281) ? 639:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1283) ? 640:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1285) ? 641:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1287) ? 642:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1289) ? 643:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1291) ? 644:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1293) ? 645:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1295) ? 646:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1297) ? 647:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1299) ? 648:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1301) ? 649:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1303) ? 650:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1305) ? 651:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1307) ? 652:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1309) ? 653:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1311) ? 654:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1313) ? 655:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1315) ? 656:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1317) ? 657:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1319) ? 658:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1321) ? 659:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1323) ? 660:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1325) ? 661:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1327) ? 662:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1329) ? 663:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1331) ? 664:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1333) ? 665:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1335) ? 666:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1337) ? 667:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1339) ? 668:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1341) ? 669:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1343) ? 670:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1345) ? 671:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1347) ? 672:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1349) ? 673:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1351) ? 674:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1353) ? 675:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1355) ? 676:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1357) ? 677:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1359) ? 678:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1361) ? 679:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1363) ? 680:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1365) ? 681:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1367) ? 682:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1369) ? 683:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1371) ? 684:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1373) ? 685:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1375) ? 686:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1377) ? 687:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1379) ? 688:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1381) ? 689:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1383) ? 690:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1385) ? 691:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1387) ? 692:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1389) ? 693:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1391) ? 694:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1393) ? 695:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1395) ? 696:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1397) ? 697:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1399) ? 698:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1401) ? 699:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1403) ? 700:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1405) ? 701:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1407) ? 702:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1409) ? 703:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1411) ? 704:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1413) ? 705:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1415) ? 706:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1417) ? 707:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1419) ? 708:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1421) ? 709:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1423) ? 710:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1425) ? 711:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1427) ? 712:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1429) ? 713:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1431) ? 714:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1433) ? 715:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1435) ? 716:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1437) ? 717:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1439) ? 718:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1441) ? 719:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1443) ? 720:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1445) ? 721:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1447) ? 722:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1449) ? 723:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1451) ? 724:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1453) ? 725:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1455) ? 726:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1457) ? 727:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1459) ? 728:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1461) ? 729:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1463) ? 730:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1465) ? 731:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1467) ? 732:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1469) ? 733:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1471) ? 734:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1473) ? 735:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1475) ? 736:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1477) ? 737:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1479) ? 738:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1481) ? 739:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1483) ? 740:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1485) ? 741:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1487) ? 742:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1489) ? 743:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1491) ? 744:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1493) ? 745:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1495) ? 746:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1497) ? 747:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1499) ? 748:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1501) ? 749:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1503) ? 750:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1505) ? 751:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1507) ? 752:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1509) ? 753:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1511) ? 754:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1513) ? 755:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1515) ? 756:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1517) ? 757:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1519) ? 758:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1521) ? 759:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1523) ? 760:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1525) ? 761:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1527) ? 762:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1529) ? 763:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1531) ? 764:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1533) ? 765:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1535) ? 766:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1537) ? 767:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1539) ? 768:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1541) ? 769:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1543) ? 770:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1545) ? 771:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1547) ? 772:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1549) ? 773:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1551) ? 774:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1553) ? 775:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1555) ? 776:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1557) ? 777:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1559) ? 778:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1561) ? 779:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1563) ? 780:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1565) ? 781:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1567) ? 782:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1569) ? 783:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1571) ? 784:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1573) ? 785:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1575) ? 786:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1577) ? 787:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1579) ? 788:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1581) ? 789:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1583) ? 790:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1585) ? 791:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1587) ? 792:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1589) ? 793:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1591) ? 794:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1593) ? 795:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1595) ? 796:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1597) ? 797:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1599) ? 798:
		       /**/
		       (r_state == zStateColumn) & (r_counter == 1601) ? 799:
		       /**/
		       0;
   assign i_raddr_beta=/**/
		       (r_counter == 0) ? 1:
		       /**/
		       (r_counter == 1) ? 2:
		       /**/
		       (r_counter == 2) ? 3:
		       /**/
		       (r_counter == 3) ? 0:
		       /**/
		       (r_counter == 4) ? 2:
		       /**/
		       (r_counter == 5) ? 3:
		       /**/
		       (r_counter == 6) ? 0:
		       /**/
		       (r_counter == 7) ? 1:
		       /**/
		       (r_counter == 8) ? 3:
		       /**/
		       (r_counter == 9) ? 0:
		       /**/
		       (r_counter == 10) ? 1:
		       /**/
		       (r_counter == 11) ? 2:
		       /**/
		       (r_counter == 12) ? 5:
		       /**/
		       (r_counter == 13) ? 6:
		       /**/
		       (r_counter == 14) ? 7:
		       /**/
		       (r_counter == 15) ? 4:
		       /**/
		       (r_counter == 16) ? 6:
		       /**/
		       (r_counter == 17) ? 7:
		       /**/
		       (r_counter == 18) ? 4:
		       /**/
		       (r_counter == 19) ? 5:
		       /**/
		       (r_counter == 20) ? 7:
		       /**/
		       (r_counter == 21) ? 4:
		       /**/
		       (r_counter == 22) ? 5:
		       /**/
		       (r_counter == 23) ? 6:
		       /**/
		       (r_counter == 24) ? 9:
		       /**/
		       (r_counter == 25) ? 10:
		       /**/
		       (r_counter == 26) ? 11:
		       /**/
		       (r_counter == 27) ? 8:
		       /**/
		       (r_counter == 28) ? 10:
		       /**/
		       (r_counter == 29) ? 11:
		       /**/
		       (r_counter == 30) ? 8:
		       /**/
		       (r_counter == 31) ? 9:
		       /**/
		       (r_counter == 32) ? 11:
		       /**/
		       (r_counter == 33) ? 8:
		       /**/
		       (r_counter == 34) ? 9:
		       /**/
		       (r_counter == 35) ? 10:
		       /**/
		       (r_counter == 36) ? 13:
		       /**/
		       (r_counter == 37) ? 14:
		       /**/
		       (r_counter == 38) ? 15:
		       /**/
		       (r_counter == 39) ? 12:
		       /**/
		       (r_counter == 40) ? 14:
		       /**/
		       (r_counter == 41) ? 15:
		       /**/
		       (r_counter == 42) ? 12:
		       /**/
		       (r_counter == 43) ? 13:
		       /**/
		       (r_counter == 44) ? 15:
		       /**/
		       (r_counter == 45) ? 12:
		       /**/
		       (r_counter == 46) ? 13:
		       /**/
		       (r_counter == 47) ? 14:
		       /**/
		       (r_counter == 48) ? 17:
		       /**/
		       (r_counter == 49) ? 18:
		       /**/
		       (r_counter == 50) ? 19:
		       /**/
		       (r_counter == 51) ? 16:
		       /**/
		       (r_counter == 52) ? 18:
		       /**/
		       (r_counter == 53) ? 19:
		       /**/
		       (r_counter == 54) ? 16:
		       /**/
		       (r_counter == 55) ? 17:
		       /**/
		       (r_counter == 56) ? 19:
		       /**/
		       (r_counter == 57) ? 16:
		       /**/
		       (r_counter == 58) ? 17:
		       /**/
		       (r_counter == 59) ? 18:
		       /**/
		       (r_counter == 60) ? 21:
		       /**/
		       (r_counter == 61) ? 22:
		       /**/
		       (r_counter == 62) ? 23:
		       /**/
		       (r_counter == 63) ? 20:
		       /**/
		       (r_counter == 64) ? 22:
		       /**/
		       (r_counter == 65) ? 23:
		       /**/
		       (r_counter == 66) ? 20:
		       /**/
		       (r_counter == 67) ? 21:
		       /**/
		       (r_counter == 68) ? 23:
		       /**/
		       (r_counter == 69) ? 20:
		       /**/
		       (r_counter == 70) ? 21:
		       /**/
		       (r_counter == 71) ? 22:
		       /**/
		       (r_counter == 72) ? 25:
		       /**/
		       (r_counter == 73) ? 26:
		       /**/
		       (r_counter == 74) ? 27:
		       /**/
		       (r_counter == 75) ? 24:
		       /**/
		       (r_counter == 76) ? 26:
		       /**/
		       (r_counter == 77) ? 27:
		       /**/
		       (r_counter == 78) ? 24:
		       /**/
		       (r_counter == 79) ? 25:
		       /**/
		       (r_counter == 80) ? 27:
		       /**/
		       (r_counter == 81) ? 24:
		       /**/
		       (r_counter == 82) ? 25:
		       /**/
		       (r_counter == 83) ? 26:
		       /**/
		       (r_counter == 84) ? 29:
		       /**/
		       (r_counter == 85) ? 30:
		       /**/
		       (r_counter == 86) ? 31:
		       /**/
		       (r_counter == 87) ? 28:
		       /**/
		       (r_counter == 88) ? 30:
		       /**/
		       (r_counter == 89) ? 31:
		       /**/
		       (r_counter == 90) ? 28:
		       /**/
		       (r_counter == 91) ? 29:
		       /**/
		       (r_counter == 92) ? 31:
		       /**/
		       (r_counter == 93) ? 28:
		       /**/
		       (r_counter == 94) ? 29:
		       /**/
		       (r_counter == 95) ? 30:
		       /**/
		       (r_counter == 96) ? 33:
		       /**/
		       (r_counter == 97) ? 34:
		       /**/
		       (r_counter == 98) ? 35:
		       /**/
		       (r_counter == 99) ? 32:
		       /**/
		       (r_counter == 100) ? 34:
		       /**/
		       (r_counter == 101) ? 35:
		       /**/
		       (r_counter == 102) ? 32:
		       /**/
		       (r_counter == 103) ? 33:
		       /**/
		       (r_counter == 104) ? 35:
		       /**/
		       (r_counter == 105) ? 32:
		       /**/
		       (r_counter == 106) ? 33:
		       /**/
		       (r_counter == 107) ? 34:
		       /**/
		       (r_counter == 108) ? 37:
		       /**/
		       (r_counter == 109) ? 38:
		       /**/
		       (r_counter == 110) ? 39:
		       /**/
		       (r_counter == 111) ? 36:
		       /**/
		       (r_counter == 112) ? 38:
		       /**/
		       (r_counter == 113) ? 39:
		       /**/
		       (r_counter == 114) ? 36:
		       /**/
		       (r_counter == 115) ? 37:
		       /**/
		       (r_counter == 116) ? 39:
		       /**/
		       (r_counter == 117) ? 36:
		       /**/
		       (r_counter == 118) ? 37:
		       /**/
		       (r_counter == 119) ? 38:
		       /**/
		       (r_counter == 120) ? 41:
		       /**/
		       (r_counter == 121) ? 42:
		       /**/
		       (r_counter == 122) ? 43:
		       /**/
		       (r_counter == 123) ? 40:
		       /**/
		       (r_counter == 124) ? 42:
		       /**/
		       (r_counter == 125) ? 43:
		       /**/
		       (r_counter == 126) ? 40:
		       /**/
		       (r_counter == 127) ? 41:
		       /**/
		       (r_counter == 128) ? 43:
		       /**/
		       (r_counter == 129) ? 40:
		       /**/
		       (r_counter == 130) ? 41:
		       /**/
		       (r_counter == 131) ? 42:
		       /**/
		       (r_counter == 132) ? 45:
		       /**/
		       (r_counter == 133) ? 46:
		       /**/
		       (r_counter == 134) ? 47:
		       /**/
		       (r_counter == 135) ? 44:
		       /**/
		       (r_counter == 136) ? 46:
		       /**/
		       (r_counter == 137) ? 47:
		       /**/
		       (r_counter == 138) ? 44:
		       /**/
		       (r_counter == 139) ? 45:
		       /**/
		       (r_counter == 140) ? 47:
		       /**/
		       (r_counter == 141) ? 44:
		       /**/
		       (r_counter == 142) ? 45:
		       /**/
		       (r_counter == 143) ? 46:
		       /**/
		       (r_counter == 144) ? 49:
		       /**/
		       (r_counter == 145) ? 50:
		       /**/
		       (r_counter == 146) ? 51:
		       /**/
		       (r_counter == 147) ? 48:
		       /**/
		       (r_counter == 148) ? 50:
		       /**/
		       (r_counter == 149) ? 51:
		       /**/
		       (r_counter == 150) ? 48:
		       /**/
		       (r_counter == 151) ? 49:
		       /**/
		       (r_counter == 152) ? 51:
		       /**/
		       (r_counter == 153) ? 48:
		       /**/
		       (r_counter == 154) ? 49:
		       /**/
		       (r_counter == 155) ? 50:
		       /**/
		       (r_counter == 156) ? 53:
		       /**/
		       (r_counter == 157) ? 54:
		       /**/
		       (r_counter == 158) ? 55:
		       /**/
		       (r_counter == 159) ? 52:
		       /**/
		       (r_counter == 160) ? 54:
		       /**/
		       (r_counter == 161) ? 55:
		       /**/
		       (r_counter == 162) ? 52:
		       /**/
		       (r_counter == 163) ? 53:
		       /**/
		       (r_counter == 164) ? 55:
		       /**/
		       (r_counter == 165) ? 52:
		       /**/
		       (r_counter == 166) ? 53:
		       /**/
		       (r_counter == 167) ? 54:
		       /**/
		       (r_counter == 168) ? 57:
		       /**/
		       (r_counter == 169) ? 58:
		       /**/
		       (r_counter == 170) ? 59:
		       /**/
		       (r_counter == 171) ? 56:
		       /**/
		       (r_counter == 172) ? 58:
		       /**/
		       (r_counter == 173) ? 59:
		       /**/
		       (r_counter == 174) ? 56:
		       /**/
		       (r_counter == 175) ? 57:
		       /**/
		       (r_counter == 176) ? 59:
		       /**/
		       (r_counter == 177) ? 56:
		       /**/
		       (r_counter == 178) ? 57:
		       /**/
		       (r_counter == 179) ? 58:
		       /**/
		       (r_counter == 180) ? 61:
		       /**/
		       (r_counter == 181) ? 62:
		       /**/
		       (r_counter == 182) ? 63:
		       /**/
		       (r_counter == 183) ? 60:
		       /**/
		       (r_counter == 184) ? 62:
		       /**/
		       (r_counter == 185) ? 63:
		       /**/
		       (r_counter == 186) ? 60:
		       /**/
		       (r_counter == 187) ? 61:
		       /**/
		       (r_counter == 188) ? 63:
		       /**/
		       (r_counter == 189) ? 60:
		       /**/
		       (r_counter == 190) ? 61:
		       /**/
		       (r_counter == 191) ? 62:
		       /**/
		       (r_counter == 192) ? 65:
		       /**/
		       (r_counter == 193) ? 66:
		       /**/
		       (r_counter == 194) ? 67:
		       /**/
		       (r_counter == 195) ? 64:
		       /**/
		       (r_counter == 196) ? 66:
		       /**/
		       (r_counter == 197) ? 67:
		       /**/
		       (r_counter == 198) ? 64:
		       /**/
		       (r_counter == 199) ? 65:
		       /**/
		       (r_counter == 200) ? 67:
		       /**/
		       (r_counter == 201) ? 64:
		       /**/
		       (r_counter == 202) ? 65:
		       /**/
		       (r_counter == 203) ? 66:
		       /**/
		       (r_counter == 204) ? 69:
		       /**/
		       (r_counter == 205) ? 70:
		       /**/
		       (r_counter == 206) ? 71:
		       /**/
		       (r_counter == 207) ? 68:
		       /**/
		       (r_counter == 208) ? 70:
		       /**/
		       (r_counter == 209) ? 71:
		       /**/
		       (r_counter == 210) ? 68:
		       /**/
		       (r_counter == 211) ? 69:
		       /**/
		       (r_counter == 212) ? 71:
		       /**/
		       (r_counter == 213) ? 68:
		       /**/
		       (r_counter == 214) ? 69:
		       /**/
		       (r_counter == 215) ? 70:
		       /**/
		       (r_counter == 216) ? 73:
		       /**/
		       (r_counter == 217) ? 74:
		       /**/
		       (r_counter == 218) ? 75:
		       /**/
		       (r_counter == 219) ? 72:
		       /**/
		       (r_counter == 220) ? 74:
		       /**/
		       (r_counter == 221) ? 75:
		       /**/
		       (r_counter == 222) ? 72:
		       /**/
		       (r_counter == 223) ? 73:
		       /**/
		       (r_counter == 224) ? 75:
		       /**/
		       (r_counter == 225) ? 72:
		       /**/
		       (r_counter == 226) ? 73:
		       /**/
		       (r_counter == 227) ? 74:
		       /**/
		       (r_counter == 228) ? 77:
		       /**/
		       (r_counter == 229) ? 78:
		       /**/
		       (r_counter == 230) ? 79:
		       /**/
		       (r_counter == 231) ? 76:
		       /**/
		       (r_counter == 232) ? 78:
		       /**/
		       (r_counter == 233) ? 79:
		       /**/
		       (r_counter == 234) ? 76:
		       /**/
		       (r_counter == 235) ? 77:
		       /**/
		       (r_counter == 236) ? 79:
		       /**/
		       (r_counter == 237) ? 76:
		       /**/
		       (r_counter == 238) ? 77:
		       /**/
		       (r_counter == 239) ? 78:
		       /**/
		       (r_counter == 240) ? 81:
		       /**/
		       (r_counter == 241) ? 82:
		       /**/
		       (r_counter == 242) ? 83:
		       /**/
		       (r_counter == 243) ? 80:
		       /**/
		       (r_counter == 244) ? 82:
		       /**/
		       (r_counter == 245) ? 83:
		       /**/
		       (r_counter == 246) ? 80:
		       /**/
		       (r_counter == 247) ? 81:
		       /**/
		       (r_counter == 248) ? 83:
		       /**/
		       (r_counter == 249) ? 80:
		       /**/
		       (r_counter == 250) ? 81:
		       /**/
		       (r_counter == 251) ? 82:
		       /**/
		       (r_counter == 252) ? 85:
		       /**/
		       (r_counter == 253) ? 86:
		       /**/
		       (r_counter == 254) ? 87:
		       /**/
		       (r_counter == 255) ? 84:
		       /**/
		       (r_counter == 256) ? 86:
		       /**/
		       (r_counter == 257) ? 87:
		       /**/
		       (r_counter == 258) ? 84:
		       /**/
		       (r_counter == 259) ? 85:
		       /**/
		       (r_counter == 260) ? 87:
		       /**/
		       (r_counter == 261) ? 84:
		       /**/
		       (r_counter == 262) ? 85:
		       /**/
		       (r_counter == 263) ? 86:
		       /**/
		       (r_counter == 264) ? 89:
		       /**/
		       (r_counter == 265) ? 90:
		       /**/
		       (r_counter == 266) ? 91:
		       /**/
		       (r_counter == 267) ? 88:
		       /**/
		       (r_counter == 268) ? 90:
		       /**/
		       (r_counter == 269) ? 91:
		       /**/
		       (r_counter == 270) ? 88:
		       /**/
		       (r_counter == 271) ? 89:
		       /**/
		       (r_counter == 272) ? 91:
		       /**/
		       (r_counter == 273) ? 88:
		       /**/
		       (r_counter == 274) ? 89:
		       /**/
		       (r_counter == 275) ? 90:
		       /**/
		       (r_counter == 276) ? 93:
		       /**/
		       (r_counter == 277) ? 94:
		       /**/
		       (r_counter == 278) ? 95:
		       /**/
		       (r_counter == 279) ? 92:
		       /**/
		       (r_counter == 280) ? 94:
		       /**/
		       (r_counter == 281) ? 95:
		       /**/
		       (r_counter == 282) ? 92:
		       /**/
		       (r_counter == 283) ? 93:
		       /**/
		       (r_counter == 284) ? 95:
		       /**/
		       (r_counter == 285) ? 92:
		       /**/
		       (r_counter == 286) ? 93:
		       /**/
		       (r_counter == 287) ? 94:
		       /**/
		       (r_counter == 288) ? 97:
		       /**/
		       (r_counter == 289) ? 98:
		       /**/
		       (r_counter == 290) ? 99:
		       /**/
		       (r_counter == 291) ? 96:
		       /**/
		       (r_counter == 292) ? 98:
		       /**/
		       (r_counter == 293) ? 99:
		       /**/
		       (r_counter == 294) ? 96:
		       /**/
		       (r_counter == 295) ? 97:
		       /**/
		       (r_counter == 296) ? 99:
		       /**/
		       (r_counter == 297) ? 96:
		       /**/
		       (r_counter == 298) ? 97:
		       /**/
		       (r_counter == 299) ? 98:
		       /**/
		       (r_counter == 300) ? 101:
		       /**/
		       (r_counter == 301) ? 102:
		       /**/
		       (r_counter == 302) ? 103:
		       /**/
		       (r_counter == 303) ? 100:
		       /**/
		       (r_counter == 304) ? 102:
		       /**/
		       (r_counter == 305) ? 103:
		       /**/
		       (r_counter == 306) ? 100:
		       /**/
		       (r_counter == 307) ? 101:
		       /**/
		       (r_counter == 308) ? 103:
		       /**/
		       (r_counter == 309) ? 100:
		       /**/
		       (r_counter == 310) ? 101:
		       /**/
		       (r_counter == 311) ? 102:
		       /**/
		       (r_counter == 312) ? 105:
		       /**/
		       (r_counter == 313) ? 106:
		       /**/
		       (r_counter == 314) ? 107:
		       /**/
		       (r_counter == 315) ? 104:
		       /**/
		       (r_counter == 316) ? 106:
		       /**/
		       (r_counter == 317) ? 107:
		       /**/
		       (r_counter == 318) ? 104:
		       /**/
		       (r_counter == 319) ? 105:
		       /**/
		       (r_counter == 320) ? 107:
		       /**/
		       (r_counter == 321) ? 104:
		       /**/
		       (r_counter == 322) ? 105:
		       /**/
		       (r_counter == 323) ? 106:
		       /**/
		       (r_counter == 324) ? 109:
		       /**/
		       (r_counter == 325) ? 110:
		       /**/
		       (r_counter == 326) ? 111:
		       /**/
		       (r_counter == 327) ? 108:
		       /**/
		       (r_counter == 328) ? 110:
		       /**/
		       (r_counter == 329) ? 111:
		       /**/
		       (r_counter == 330) ? 108:
		       /**/
		       (r_counter == 331) ? 109:
		       /**/
		       (r_counter == 332) ? 111:
		       /**/
		       (r_counter == 333) ? 108:
		       /**/
		       (r_counter == 334) ? 109:
		       /**/
		       (r_counter == 335) ? 110:
		       /**/
		       (r_counter == 336) ? 113:
		       /**/
		       (r_counter == 337) ? 114:
		       /**/
		       (r_counter == 338) ? 115:
		       /**/
		       (r_counter == 339) ? 112:
		       /**/
		       (r_counter == 340) ? 114:
		       /**/
		       (r_counter == 341) ? 115:
		       /**/
		       (r_counter == 342) ? 112:
		       /**/
		       (r_counter == 343) ? 113:
		       /**/
		       (r_counter == 344) ? 115:
		       /**/
		       (r_counter == 345) ? 112:
		       /**/
		       (r_counter == 346) ? 113:
		       /**/
		       (r_counter == 347) ? 114:
		       /**/
		       (r_counter == 348) ? 117:
		       /**/
		       (r_counter == 349) ? 118:
		       /**/
		       (r_counter == 350) ? 119:
		       /**/
		       (r_counter == 351) ? 116:
		       /**/
		       (r_counter == 352) ? 118:
		       /**/
		       (r_counter == 353) ? 119:
		       /**/
		       (r_counter == 354) ? 116:
		       /**/
		       (r_counter == 355) ? 117:
		       /**/
		       (r_counter == 356) ? 119:
		       /**/
		       (r_counter == 357) ? 116:
		       /**/
		       (r_counter == 358) ? 117:
		       /**/
		       (r_counter == 359) ? 118:
		       /**/
		       (r_counter == 360) ? 121:
		       /**/
		       (r_counter == 361) ? 122:
		       /**/
		       (r_counter == 362) ? 123:
		       /**/
		       (r_counter == 363) ? 120:
		       /**/
		       (r_counter == 364) ? 122:
		       /**/
		       (r_counter == 365) ? 123:
		       /**/
		       (r_counter == 366) ? 120:
		       /**/
		       (r_counter == 367) ? 121:
		       /**/
		       (r_counter == 368) ? 123:
		       /**/
		       (r_counter == 369) ? 120:
		       /**/
		       (r_counter == 370) ? 121:
		       /**/
		       (r_counter == 371) ? 122:
		       /**/
		       (r_counter == 372) ? 125:
		       /**/
		       (r_counter == 373) ? 126:
		       /**/
		       (r_counter == 374) ? 127:
		       /**/
		       (r_counter == 375) ? 124:
		       /**/
		       (r_counter == 376) ? 126:
		       /**/
		       (r_counter == 377) ? 127:
		       /**/
		       (r_counter == 378) ? 124:
		       /**/
		       (r_counter == 379) ? 125:
		       /**/
		       (r_counter == 380) ? 127:
		       /**/
		       (r_counter == 381) ? 124:
		       /**/
		       (r_counter == 382) ? 125:
		       /**/
		       (r_counter == 383) ? 126:
		       /**/
		       (r_counter == 384) ? 129:
		       /**/
		       (r_counter == 385) ? 130:
		       /**/
		       (r_counter == 386) ? 131:
		       /**/
		       (r_counter == 387) ? 128:
		       /**/
		       (r_counter == 388) ? 130:
		       /**/
		       (r_counter == 389) ? 131:
		       /**/
		       (r_counter == 390) ? 128:
		       /**/
		       (r_counter == 391) ? 129:
		       /**/
		       (r_counter == 392) ? 131:
		       /**/
		       (r_counter == 393) ? 128:
		       /**/
		       (r_counter == 394) ? 129:
		       /**/
		       (r_counter == 395) ? 130:
		       /**/
		       (r_counter == 396) ? 133:
		       /**/
		       (r_counter == 397) ? 134:
		       /**/
		       (r_counter == 398) ? 135:
		       /**/
		       (r_counter == 399) ? 132:
		       /**/
		       (r_counter == 400) ? 134:
		       /**/
		       (r_counter == 401) ? 135:
		       /**/
		       (r_counter == 402) ? 132:
		       /**/
		       (r_counter == 403) ? 133:
		       /**/
		       (r_counter == 404) ? 135:
		       /**/
		       (r_counter == 405) ? 132:
		       /**/
		       (r_counter == 406) ? 133:
		       /**/
		       (r_counter == 407) ? 134:
		       /**/
		       (r_counter == 408) ? 137:
		       /**/
		       (r_counter == 409) ? 138:
		       /**/
		       (r_counter == 410) ? 139:
		       /**/
		       (r_counter == 411) ? 136:
		       /**/
		       (r_counter == 412) ? 138:
		       /**/
		       (r_counter == 413) ? 139:
		       /**/
		       (r_counter == 414) ? 136:
		       /**/
		       (r_counter == 415) ? 137:
		       /**/
		       (r_counter == 416) ? 139:
		       /**/
		       (r_counter == 417) ? 136:
		       /**/
		       (r_counter == 418) ? 137:
		       /**/
		       (r_counter == 419) ? 138:
		       /**/
		       (r_counter == 420) ? 141:
		       /**/
		       (r_counter == 421) ? 142:
		       /**/
		       (r_counter == 422) ? 143:
		       /**/
		       (r_counter == 423) ? 140:
		       /**/
		       (r_counter == 424) ? 142:
		       /**/
		       (r_counter == 425) ? 143:
		       /**/
		       (r_counter == 426) ? 140:
		       /**/
		       (r_counter == 427) ? 141:
		       /**/
		       (r_counter == 428) ? 143:
		       /**/
		       (r_counter == 429) ? 140:
		       /**/
		       (r_counter == 430) ? 141:
		       /**/
		       (r_counter == 431) ? 142:
		       /**/
		       (r_counter == 432) ? 145:
		       /**/
		       (r_counter == 433) ? 146:
		       /**/
		       (r_counter == 434) ? 147:
		       /**/
		       (r_counter == 435) ? 144:
		       /**/
		       (r_counter == 436) ? 146:
		       /**/
		       (r_counter == 437) ? 147:
		       /**/
		       (r_counter == 438) ? 144:
		       /**/
		       (r_counter == 439) ? 145:
		       /**/
		       (r_counter == 440) ? 147:
		       /**/
		       (r_counter == 441) ? 144:
		       /**/
		       (r_counter == 442) ? 145:
		       /**/
		       (r_counter == 443) ? 146:
		       /**/
		       (r_counter == 444) ? 149:
		       /**/
		       (r_counter == 445) ? 150:
		       /**/
		       (r_counter == 446) ? 151:
		       /**/
		       (r_counter == 447) ? 148:
		       /**/
		       (r_counter == 448) ? 150:
		       /**/
		       (r_counter == 449) ? 151:
		       /**/
		       (r_counter == 450) ? 148:
		       /**/
		       (r_counter == 451) ? 149:
		       /**/
		       (r_counter == 452) ? 151:
		       /**/
		       (r_counter == 453) ? 148:
		       /**/
		       (r_counter == 454) ? 149:
		       /**/
		       (r_counter == 455) ? 150:
		       /**/
		       (r_counter == 456) ? 153:
		       /**/
		       (r_counter == 457) ? 154:
		       /**/
		       (r_counter == 458) ? 155:
		       /**/
		       (r_counter == 459) ? 152:
		       /**/
		       (r_counter == 460) ? 154:
		       /**/
		       (r_counter == 461) ? 155:
		       /**/
		       (r_counter == 462) ? 152:
		       /**/
		       (r_counter == 463) ? 153:
		       /**/
		       (r_counter == 464) ? 155:
		       /**/
		       (r_counter == 465) ? 152:
		       /**/
		       (r_counter == 466) ? 153:
		       /**/
		       (r_counter == 467) ? 154:
		       /**/
		       (r_counter == 468) ? 157:
		       /**/
		       (r_counter == 469) ? 158:
		       /**/
		       (r_counter == 470) ? 159:
		       /**/
		       (r_counter == 471) ? 156:
		       /**/
		       (r_counter == 472) ? 158:
		       /**/
		       (r_counter == 473) ? 159:
		       /**/
		       (r_counter == 474) ? 156:
		       /**/
		       (r_counter == 475) ? 157:
		       /**/
		       (r_counter == 476) ? 159:
		       /**/
		       (r_counter == 477) ? 156:
		       /**/
		       (r_counter == 478) ? 157:
		       /**/
		       (r_counter == 479) ? 158:
		       /**/
		       (r_counter == 480) ? 161:
		       /**/
		       (r_counter == 481) ? 162:
		       /**/
		       (r_counter == 482) ? 163:
		       /**/
		       (r_counter == 483) ? 160:
		       /**/
		       (r_counter == 484) ? 162:
		       /**/
		       (r_counter == 485) ? 163:
		       /**/
		       (r_counter == 486) ? 160:
		       /**/
		       (r_counter == 487) ? 161:
		       /**/
		       (r_counter == 488) ? 163:
		       /**/
		       (r_counter == 489) ? 160:
		       /**/
		       (r_counter == 490) ? 161:
		       /**/
		       (r_counter == 491) ? 162:
		       /**/
		       (r_counter == 492) ? 165:
		       /**/
		       (r_counter == 493) ? 166:
		       /**/
		       (r_counter == 494) ? 167:
		       /**/
		       (r_counter == 495) ? 164:
		       /**/
		       (r_counter == 496) ? 166:
		       /**/
		       (r_counter == 497) ? 167:
		       /**/
		       (r_counter == 498) ? 164:
		       /**/
		       (r_counter == 499) ? 165:
		       /**/
		       (r_counter == 500) ? 167:
		       /**/
		       (r_counter == 501) ? 164:
		       /**/
		       (r_counter == 502) ? 165:
		       /**/
		       (r_counter == 503) ? 166:
		       /**/
		       (r_counter == 504) ? 169:
		       /**/
		       (r_counter == 505) ? 170:
		       /**/
		       (r_counter == 506) ? 171:
		       /**/
		       (r_counter == 507) ? 168:
		       /**/
		       (r_counter == 508) ? 170:
		       /**/
		       (r_counter == 509) ? 171:
		       /**/
		       (r_counter == 510) ? 168:
		       /**/
		       (r_counter == 511) ? 169:
		       /**/
		       (r_counter == 512) ? 171:
		       /**/
		       (r_counter == 513) ? 168:
		       /**/
		       (r_counter == 514) ? 169:
		       /**/
		       (r_counter == 515) ? 170:
		       /**/
		       (r_counter == 516) ? 173:
		       /**/
		       (r_counter == 517) ? 174:
		       /**/
		       (r_counter == 518) ? 175:
		       /**/
		       (r_counter == 519) ? 172:
		       /**/
		       (r_counter == 520) ? 174:
		       /**/
		       (r_counter == 521) ? 175:
		       /**/
		       (r_counter == 522) ? 172:
		       /**/
		       (r_counter == 523) ? 173:
		       /**/
		       (r_counter == 524) ? 175:
		       /**/
		       (r_counter == 525) ? 172:
		       /**/
		       (r_counter == 526) ? 173:
		       /**/
		       (r_counter == 527) ? 174:
		       /**/
		       (r_counter == 528) ? 177:
		       /**/
		       (r_counter == 529) ? 178:
		       /**/
		       (r_counter == 530) ? 179:
		       /**/
		       (r_counter == 531) ? 176:
		       /**/
		       (r_counter == 532) ? 178:
		       /**/
		       (r_counter == 533) ? 179:
		       /**/
		       (r_counter == 534) ? 176:
		       /**/
		       (r_counter == 535) ? 177:
		       /**/
		       (r_counter == 536) ? 179:
		       /**/
		       (r_counter == 537) ? 176:
		       /**/
		       (r_counter == 538) ? 177:
		       /**/
		       (r_counter == 539) ? 178:
		       /**/
		       (r_counter == 540) ? 181:
		       /**/
		       (r_counter == 541) ? 182:
		       /**/
		       (r_counter == 542) ? 183:
		       /**/
		       (r_counter == 543) ? 180:
		       /**/
		       (r_counter == 544) ? 182:
		       /**/
		       (r_counter == 545) ? 183:
		       /**/
		       (r_counter == 546) ? 180:
		       /**/
		       (r_counter == 547) ? 181:
		       /**/
		       (r_counter == 548) ? 183:
		       /**/
		       (r_counter == 549) ? 180:
		       /**/
		       (r_counter == 550) ? 181:
		       /**/
		       (r_counter == 551) ? 182:
		       /**/
		       (r_counter == 552) ? 185:
		       /**/
		       (r_counter == 553) ? 186:
		       /**/
		       (r_counter == 554) ? 187:
		       /**/
		       (r_counter == 555) ? 184:
		       /**/
		       (r_counter == 556) ? 186:
		       /**/
		       (r_counter == 557) ? 187:
		       /**/
		       (r_counter == 558) ? 184:
		       /**/
		       (r_counter == 559) ? 185:
		       /**/
		       (r_counter == 560) ? 187:
		       /**/
		       (r_counter == 561) ? 184:
		       /**/
		       (r_counter == 562) ? 185:
		       /**/
		       (r_counter == 563) ? 186:
		       /**/
		       (r_counter == 564) ? 189:
		       /**/
		       (r_counter == 565) ? 190:
		       /**/
		       (r_counter == 566) ? 191:
		       /**/
		       (r_counter == 567) ? 188:
		       /**/
		       (r_counter == 568) ? 190:
		       /**/
		       (r_counter == 569) ? 191:
		       /**/
		       (r_counter == 570) ? 188:
		       /**/
		       (r_counter == 571) ? 189:
		       /**/
		       (r_counter == 572) ? 191:
		       /**/
		       (r_counter == 573) ? 188:
		       /**/
		       (r_counter == 574) ? 189:
		       /**/
		       (r_counter == 575) ? 190:
		       /**/
		       (r_counter == 576) ? 193:
		       /**/
		       (r_counter == 577) ? 194:
		       /**/
		       (r_counter == 578) ? 195:
		       /**/
		       (r_counter == 579) ? 192:
		       /**/
		       (r_counter == 580) ? 194:
		       /**/
		       (r_counter == 581) ? 195:
		       /**/
		       (r_counter == 582) ? 192:
		       /**/
		       (r_counter == 583) ? 193:
		       /**/
		       (r_counter == 584) ? 195:
		       /**/
		       (r_counter == 585) ? 192:
		       /**/
		       (r_counter == 586) ? 193:
		       /**/
		       (r_counter == 587) ? 194:
		       /**/
		       (r_counter == 588) ? 197:
		       /**/
		       (r_counter == 589) ? 198:
		       /**/
		       (r_counter == 590) ? 199:
		       /**/
		       (r_counter == 591) ? 196:
		       /**/
		       (r_counter == 592) ? 198:
		       /**/
		       (r_counter == 593) ? 199:
		       /**/
		       (r_counter == 594) ? 196:
		       /**/
		       (r_counter == 595) ? 197:
		       /**/
		       (r_counter == 596) ? 199:
		       /**/
		       (r_counter == 597) ? 196:
		       /**/
		       (r_counter == 598) ? 197:
		       /**/
		       (r_counter == 599) ? 198:
		       /**/
		       (r_counter == 600) ? 201:
		       /**/
		       (r_counter == 601) ? 202:
		       /**/
		       (r_counter == 602) ? 203:
		       /**/
		       (r_counter == 603) ? 200:
		       /**/
		       (r_counter == 604) ? 202:
		       /**/
		       (r_counter == 605) ? 203:
		       /**/
		       (r_counter == 606) ? 200:
		       /**/
		       (r_counter == 607) ? 201:
		       /**/
		       (r_counter == 608) ? 203:
		       /**/
		       (r_counter == 609) ? 200:
		       /**/
		       (r_counter == 610) ? 201:
		       /**/
		       (r_counter == 611) ? 202:
		       /**/
		       (r_counter == 612) ? 205:
		       /**/
		       (r_counter == 613) ? 206:
		       /**/
		       (r_counter == 614) ? 207:
		       /**/
		       (r_counter == 615) ? 204:
		       /**/
		       (r_counter == 616) ? 206:
		       /**/
		       (r_counter == 617) ? 207:
		       /**/
		       (r_counter == 618) ? 204:
		       /**/
		       (r_counter == 619) ? 205:
		       /**/
		       (r_counter == 620) ? 207:
		       /**/
		       (r_counter == 621) ? 204:
		       /**/
		       (r_counter == 622) ? 205:
		       /**/
		       (r_counter == 623) ? 206:
		       /**/
		       (r_counter == 624) ? 209:
		       /**/
		       (r_counter == 625) ? 210:
		       /**/
		       (r_counter == 626) ? 211:
		       /**/
		       (r_counter == 627) ? 208:
		       /**/
		       (r_counter == 628) ? 210:
		       /**/
		       (r_counter == 629) ? 211:
		       /**/
		       (r_counter == 630) ? 208:
		       /**/
		       (r_counter == 631) ? 209:
		       /**/
		       (r_counter == 632) ? 211:
		       /**/
		       (r_counter == 633) ? 208:
		       /**/
		       (r_counter == 634) ? 209:
		       /**/
		       (r_counter == 635) ? 210:
		       /**/
		       (r_counter == 636) ? 213:
		       /**/
		       (r_counter == 637) ? 214:
		       /**/
		       (r_counter == 638) ? 215:
		       /**/
		       (r_counter == 639) ? 212:
		       /**/
		       (r_counter == 640) ? 214:
		       /**/
		       (r_counter == 641) ? 215:
		       /**/
		       (r_counter == 642) ? 212:
		       /**/
		       (r_counter == 643) ? 213:
		       /**/
		       (r_counter == 644) ? 215:
		       /**/
		       (r_counter == 645) ? 212:
		       /**/
		       (r_counter == 646) ? 213:
		       /**/
		       (r_counter == 647) ? 214:
		       /**/
		       (r_counter == 648) ? 217:
		       /**/
		       (r_counter == 649) ? 218:
		       /**/
		       (r_counter == 650) ? 219:
		       /**/
		       (r_counter == 651) ? 216:
		       /**/
		       (r_counter == 652) ? 218:
		       /**/
		       (r_counter == 653) ? 219:
		       /**/
		       (r_counter == 654) ? 216:
		       /**/
		       (r_counter == 655) ? 217:
		       /**/
		       (r_counter == 656) ? 219:
		       /**/
		       (r_counter == 657) ? 216:
		       /**/
		       (r_counter == 658) ? 217:
		       /**/
		       (r_counter == 659) ? 218:
		       /**/
		       (r_counter == 660) ? 221:
		       /**/
		       (r_counter == 661) ? 222:
		       /**/
		       (r_counter == 662) ? 223:
		       /**/
		       (r_counter == 663) ? 220:
		       /**/
		       (r_counter == 664) ? 222:
		       /**/
		       (r_counter == 665) ? 223:
		       /**/
		       (r_counter == 666) ? 220:
		       /**/
		       (r_counter == 667) ? 221:
		       /**/
		       (r_counter == 668) ? 223:
		       /**/
		       (r_counter == 669) ? 220:
		       /**/
		       (r_counter == 670) ? 221:
		       /**/
		       (r_counter == 671) ? 222:
		       /**/
		       (r_counter == 672) ? 225:
		       /**/
		       (r_counter == 673) ? 226:
		       /**/
		       (r_counter == 674) ? 227:
		       /**/
		       (r_counter == 675) ? 224:
		       /**/
		       (r_counter == 676) ? 226:
		       /**/
		       (r_counter == 677) ? 227:
		       /**/
		       (r_counter == 678) ? 224:
		       /**/
		       (r_counter == 679) ? 225:
		       /**/
		       (r_counter == 680) ? 227:
		       /**/
		       (r_counter == 681) ? 224:
		       /**/
		       (r_counter == 682) ? 225:
		       /**/
		       (r_counter == 683) ? 226:
		       /**/
		       (r_counter == 684) ? 229:
		       /**/
		       (r_counter == 685) ? 230:
		       /**/
		       (r_counter == 686) ? 231:
		       /**/
		       (r_counter == 687) ? 228:
		       /**/
		       (r_counter == 688) ? 230:
		       /**/
		       (r_counter == 689) ? 231:
		       /**/
		       (r_counter == 690) ? 228:
		       /**/
		       (r_counter == 691) ? 229:
		       /**/
		       (r_counter == 692) ? 231:
		       /**/
		       (r_counter == 693) ? 228:
		       /**/
		       (r_counter == 694) ? 229:
		       /**/
		       (r_counter == 695) ? 230:
		       /**/
		       (r_counter == 696) ? 233:
		       /**/
		       (r_counter == 697) ? 234:
		       /**/
		       (r_counter == 698) ? 235:
		       /**/
		       (r_counter == 699) ? 232:
		       /**/
		       (r_counter == 700) ? 234:
		       /**/
		       (r_counter == 701) ? 235:
		       /**/
		       (r_counter == 702) ? 232:
		       /**/
		       (r_counter == 703) ? 233:
		       /**/
		       (r_counter == 704) ? 235:
		       /**/
		       (r_counter == 705) ? 232:
		       /**/
		       (r_counter == 706) ? 233:
		       /**/
		       (r_counter == 707) ? 234:
		       /**/
		       (r_counter == 708) ? 237:
		       /**/
		       (r_counter == 709) ? 238:
		       /**/
		       (r_counter == 710) ? 239:
		       /**/
		       (r_counter == 711) ? 236:
		       /**/
		       (r_counter == 712) ? 238:
		       /**/
		       (r_counter == 713) ? 239:
		       /**/
		       (r_counter == 714) ? 236:
		       /**/
		       (r_counter == 715) ? 237:
		       /**/
		       (r_counter == 716) ? 239:
		       /**/
		       (r_counter == 717) ? 236:
		       /**/
		       (r_counter == 718) ? 237:
		       /**/
		       (r_counter == 719) ? 238:
		       /**/
		       (r_counter == 720) ? 241:
		       /**/
		       (r_counter == 721) ? 242:
		       /**/
		       (r_counter == 722) ? 243:
		       /**/
		       (r_counter == 723) ? 240:
		       /**/
		       (r_counter == 724) ? 242:
		       /**/
		       (r_counter == 725) ? 243:
		       /**/
		       (r_counter == 726) ? 240:
		       /**/
		       (r_counter == 727) ? 241:
		       /**/
		       (r_counter == 728) ? 243:
		       /**/
		       (r_counter == 729) ? 240:
		       /**/
		       (r_counter == 730) ? 241:
		       /**/
		       (r_counter == 731) ? 242:
		       /**/
		       (r_counter == 732) ? 245:
		       /**/
		       (r_counter == 733) ? 246:
		       /**/
		       (r_counter == 734) ? 247:
		       /**/
		       (r_counter == 735) ? 244:
		       /**/
		       (r_counter == 736) ? 246:
		       /**/
		       (r_counter == 737) ? 247:
		       /**/
		       (r_counter == 738) ? 244:
		       /**/
		       (r_counter == 739) ? 245:
		       /**/
		       (r_counter == 740) ? 247:
		       /**/
		       (r_counter == 741) ? 244:
		       /**/
		       (r_counter == 742) ? 245:
		       /**/
		       (r_counter == 743) ? 246:
		       /**/
		       (r_counter == 744) ? 249:
		       /**/
		       (r_counter == 745) ? 250:
		       /**/
		       (r_counter == 746) ? 251:
		       /**/
		       (r_counter == 747) ? 248:
		       /**/
		       (r_counter == 748) ? 250:
		       /**/
		       (r_counter == 749) ? 251:
		       /**/
		       (r_counter == 750) ? 248:
		       /**/
		       (r_counter == 751) ? 249:
		       /**/
		       (r_counter == 752) ? 251:
		       /**/
		       (r_counter == 753) ? 248:
		       /**/
		       (r_counter == 754) ? 249:
		       /**/
		       (r_counter == 755) ? 250:
		       /**/
		       (r_counter == 756) ? 253:
		       /**/
		       (r_counter == 757) ? 254:
		       /**/
		       (r_counter == 758) ? 255:
		       /**/
		       (r_counter == 759) ? 252:
		       /**/
		       (r_counter == 760) ? 254:
		       /**/
		       (r_counter == 761) ? 255:
		       /**/
		       (r_counter == 762) ? 252:
		       /**/
		       (r_counter == 763) ? 253:
		       /**/
		       (r_counter == 764) ? 255:
		       /**/
		       (r_counter == 765) ? 252:
		       /**/
		       (r_counter == 766) ? 253:
		       /**/
		       (r_counter == 767) ? 254:
		       /**/
		       (r_counter == 768) ? 257:
		       /**/
		       (r_counter == 769) ? 258:
		       /**/
		       (r_counter == 770) ? 259:
		       /**/
		       (r_counter == 771) ? 256:
		       /**/
		       (r_counter == 772) ? 258:
		       /**/
		       (r_counter == 773) ? 259:
		       /**/
		       (r_counter == 774) ? 256:
		       /**/
		       (r_counter == 775) ? 257:
		       /**/
		       (r_counter == 776) ? 259:
		       /**/
		       (r_counter == 777) ? 256:
		       /**/
		       (r_counter == 778) ? 257:
		       /**/
		       (r_counter == 779) ? 258:
		       /**/
		       (r_counter == 780) ? 261:
		       /**/
		       (r_counter == 781) ? 262:
		       /**/
		       (r_counter == 782) ? 263:
		       /**/
		       (r_counter == 783) ? 260:
		       /**/
		       (r_counter == 784) ? 262:
		       /**/
		       (r_counter == 785) ? 263:
		       /**/
		       (r_counter == 786) ? 260:
		       /**/
		       (r_counter == 787) ? 261:
		       /**/
		       (r_counter == 788) ? 263:
		       /**/
		       (r_counter == 789) ? 260:
		       /**/
		       (r_counter == 790) ? 261:
		       /**/
		       (r_counter == 791) ? 262:
		       /**/
		       (r_counter == 792) ? 265:
		       /**/
		       (r_counter == 793) ? 266:
		       /**/
		       (r_counter == 794) ? 267:
		       /**/
		       (r_counter == 795) ? 264:
		       /**/
		       (r_counter == 796) ? 266:
		       /**/
		       (r_counter == 797) ? 267:
		       /**/
		       (r_counter == 798) ? 264:
		       /**/
		       (r_counter == 799) ? 265:
		       /**/
		       (r_counter == 800) ? 267:
		       /**/
		       (r_counter == 801) ? 264:
		       /**/
		       (r_counter == 802) ? 265:
		       /**/
		       (r_counter == 803) ? 266:
		       /**/
		       (r_counter == 804) ? 269:
		       /**/
		       (r_counter == 805) ? 270:
		       /**/
		       (r_counter == 806) ? 271:
		       /**/
		       (r_counter == 807) ? 268:
		       /**/
		       (r_counter == 808) ? 270:
		       /**/
		       (r_counter == 809) ? 271:
		       /**/
		       (r_counter == 810) ? 268:
		       /**/
		       (r_counter == 811) ? 269:
		       /**/
		       (r_counter == 812) ? 271:
		       /**/
		       (r_counter == 813) ? 268:
		       /**/
		       (r_counter == 814) ? 269:
		       /**/
		       (r_counter == 815) ? 270:
		       /**/
		       (r_counter == 816) ? 273:
		       /**/
		       (r_counter == 817) ? 274:
		       /**/
		       (r_counter == 818) ? 275:
		       /**/
		       (r_counter == 819) ? 272:
		       /**/
		       (r_counter == 820) ? 274:
		       /**/
		       (r_counter == 821) ? 275:
		       /**/
		       (r_counter == 822) ? 272:
		       /**/
		       (r_counter == 823) ? 273:
		       /**/
		       (r_counter == 824) ? 275:
		       /**/
		       (r_counter == 825) ? 272:
		       /**/
		       (r_counter == 826) ? 273:
		       /**/
		       (r_counter == 827) ? 274:
		       /**/
		       (r_counter == 828) ? 277:
		       /**/
		       (r_counter == 829) ? 278:
		       /**/
		       (r_counter == 830) ? 279:
		       /**/
		       (r_counter == 831) ? 276:
		       /**/
		       (r_counter == 832) ? 278:
		       /**/
		       (r_counter == 833) ? 279:
		       /**/
		       (r_counter == 834) ? 276:
		       /**/
		       (r_counter == 835) ? 277:
		       /**/
		       (r_counter == 836) ? 279:
		       /**/
		       (r_counter == 837) ? 276:
		       /**/
		       (r_counter == 838) ? 277:
		       /**/
		       (r_counter == 839) ? 278:
		       /**/
		       (r_counter == 840) ? 281:
		       /**/
		       (r_counter == 841) ? 282:
		       /**/
		       (r_counter == 842) ? 283:
		       /**/
		       (r_counter == 843) ? 280:
		       /**/
		       (r_counter == 844) ? 282:
		       /**/
		       (r_counter == 845) ? 283:
		       /**/
		       (r_counter == 846) ? 280:
		       /**/
		       (r_counter == 847) ? 281:
		       /**/
		       (r_counter == 848) ? 283:
		       /**/
		       (r_counter == 849) ? 280:
		       /**/
		       (r_counter == 850) ? 281:
		       /**/
		       (r_counter == 851) ? 282:
		       /**/
		       (r_counter == 852) ? 285:
		       /**/
		       (r_counter == 853) ? 286:
		       /**/
		       (r_counter == 854) ? 287:
		       /**/
		       (r_counter == 855) ? 284:
		       /**/
		       (r_counter == 856) ? 286:
		       /**/
		       (r_counter == 857) ? 287:
		       /**/
		       (r_counter == 858) ? 284:
		       /**/
		       (r_counter == 859) ? 285:
		       /**/
		       (r_counter == 860) ? 287:
		       /**/
		       (r_counter == 861) ? 284:
		       /**/
		       (r_counter == 862) ? 285:
		       /**/
		       (r_counter == 863) ? 286:
		       /**/
		       (r_counter == 864) ? 289:
		       /**/
		       (r_counter == 865) ? 290:
		       /**/
		       (r_counter == 866) ? 291:
		       /**/
		       (r_counter == 867) ? 288:
		       /**/
		       (r_counter == 868) ? 290:
		       /**/
		       (r_counter == 869) ? 291:
		       /**/
		       (r_counter == 870) ? 288:
		       /**/
		       (r_counter == 871) ? 289:
		       /**/
		       (r_counter == 872) ? 291:
		       /**/
		       (r_counter == 873) ? 288:
		       /**/
		       (r_counter == 874) ? 289:
		       /**/
		       (r_counter == 875) ? 290:
		       /**/
		       (r_counter == 876) ? 293:
		       /**/
		       (r_counter == 877) ? 294:
		       /**/
		       (r_counter == 878) ? 295:
		       /**/
		       (r_counter == 879) ? 292:
		       /**/
		       (r_counter == 880) ? 294:
		       /**/
		       (r_counter == 881) ? 295:
		       /**/
		       (r_counter == 882) ? 292:
		       /**/
		       (r_counter == 883) ? 293:
		       /**/
		       (r_counter == 884) ? 295:
		       /**/
		       (r_counter == 885) ? 292:
		       /**/
		       (r_counter == 886) ? 293:
		       /**/
		       (r_counter == 887) ? 294:
		       /**/
		       (r_counter == 888) ? 297:
		       /**/
		       (r_counter == 889) ? 298:
		       /**/
		       (r_counter == 890) ? 299:
		       /**/
		       (r_counter == 891) ? 296:
		       /**/
		       (r_counter == 892) ? 298:
		       /**/
		       (r_counter == 893) ? 299:
		       /**/
		       (r_counter == 894) ? 296:
		       /**/
		       (r_counter == 895) ? 297:
		       /**/
		       (r_counter == 896) ? 299:
		       /**/
		       (r_counter == 897) ? 296:
		       /**/
		       (r_counter == 898) ? 297:
		       /**/
		       (r_counter == 899) ? 298:
		       /**/
		       (r_counter == 900) ? 301:
		       /**/
		       (r_counter == 901) ? 302:
		       /**/
		       (r_counter == 902) ? 303:
		       /**/
		       (r_counter == 903) ? 300:
		       /**/
		       (r_counter == 904) ? 302:
		       /**/
		       (r_counter == 905) ? 303:
		       /**/
		       (r_counter == 906) ? 300:
		       /**/
		       (r_counter == 907) ? 301:
		       /**/
		       (r_counter == 908) ? 303:
		       /**/
		       (r_counter == 909) ? 300:
		       /**/
		       (r_counter == 910) ? 301:
		       /**/
		       (r_counter == 911) ? 302:
		       /**/
		       (r_counter == 912) ? 305:
		       /**/
		       (r_counter == 913) ? 306:
		       /**/
		       (r_counter == 914) ? 307:
		       /**/
		       (r_counter == 915) ? 304:
		       /**/
		       (r_counter == 916) ? 306:
		       /**/
		       (r_counter == 917) ? 307:
		       /**/
		       (r_counter == 918) ? 304:
		       /**/
		       (r_counter == 919) ? 305:
		       /**/
		       (r_counter == 920) ? 307:
		       /**/
		       (r_counter == 921) ? 304:
		       /**/
		       (r_counter == 922) ? 305:
		       /**/
		       (r_counter == 923) ? 306:
		       /**/
		       (r_counter == 924) ? 309:
		       /**/
		       (r_counter == 925) ? 310:
		       /**/
		       (r_counter == 926) ? 311:
		       /**/
		       (r_counter == 927) ? 308:
		       /**/
		       (r_counter == 928) ? 310:
		       /**/
		       (r_counter == 929) ? 311:
		       /**/
		       (r_counter == 930) ? 308:
		       /**/
		       (r_counter == 931) ? 309:
		       /**/
		       (r_counter == 932) ? 311:
		       /**/
		       (r_counter == 933) ? 308:
		       /**/
		       (r_counter == 934) ? 309:
		       /**/
		       (r_counter == 935) ? 310:
		       /**/
		       (r_counter == 936) ? 313:
		       /**/
		       (r_counter == 937) ? 314:
		       /**/
		       (r_counter == 938) ? 315:
		       /**/
		       (r_counter == 939) ? 312:
		       /**/
		       (r_counter == 940) ? 314:
		       /**/
		       (r_counter == 941) ? 315:
		       /**/
		       (r_counter == 942) ? 312:
		       /**/
		       (r_counter == 943) ? 313:
		       /**/
		       (r_counter == 944) ? 315:
		       /**/
		       (r_counter == 945) ? 312:
		       /**/
		       (r_counter == 946) ? 313:
		       /**/
		       (r_counter == 947) ? 314:
		       /**/
		       (r_counter == 948) ? 317:
		       /**/
		       (r_counter == 949) ? 318:
		       /**/
		       (r_counter == 950) ? 319:
		       /**/
		       (r_counter == 951) ? 316:
		       /**/
		       (r_counter == 952) ? 318:
		       /**/
		       (r_counter == 953) ? 319:
		       /**/
		       (r_counter == 954) ? 316:
		       /**/
		       (r_counter == 955) ? 317:
		       /**/
		       (r_counter == 956) ? 319:
		       /**/
		       (r_counter == 957) ? 316:
		       /**/
		       (r_counter == 958) ? 317:
		       /**/
		       (r_counter == 959) ? 318:
		       /**/
		       (r_counter == 960) ? 321:
		       /**/
		       (r_counter == 961) ? 322:
		       /**/
		       (r_counter == 962) ? 323:
		       /**/
		       (r_counter == 963) ? 320:
		       /**/
		       (r_counter == 964) ? 322:
		       /**/
		       (r_counter == 965) ? 323:
		       /**/
		       (r_counter == 966) ? 320:
		       /**/
		       (r_counter == 967) ? 321:
		       /**/
		       (r_counter == 968) ? 323:
		       /**/
		       (r_counter == 969) ? 320:
		       /**/
		       (r_counter == 970) ? 321:
		       /**/
		       (r_counter == 971) ? 322:
		       /**/
		       (r_counter == 972) ? 325:
		       /**/
		       (r_counter == 973) ? 326:
		       /**/
		       (r_counter == 974) ? 327:
		       /**/
		       (r_counter == 975) ? 324:
		       /**/
		       (r_counter == 976) ? 326:
		       /**/
		       (r_counter == 977) ? 327:
		       /**/
		       (r_counter == 978) ? 324:
		       /**/
		       (r_counter == 979) ? 325:
		       /**/
		       (r_counter == 980) ? 327:
		       /**/
		       (r_counter == 981) ? 324:
		       /**/
		       (r_counter == 982) ? 325:
		       /**/
		       (r_counter == 983) ? 326:
		       /**/
		       (r_counter == 984) ? 329:
		       /**/
		       (r_counter == 985) ? 330:
		       /**/
		       (r_counter == 986) ? 331:
		       /**/
		       (r_counter == 987) ? 328:
		       /**/
		       (r_counter == 988) ? 330:
		       /**/
		       (r_counter == 989) ? 331:
		       /**/
		       (r_counter == 990) ? 328:
		       /**/
		       (r_counter == 991) ? 329:
		       /**/
		       (r_counter == 992) ? 331:
		       /**/
		       (r_counter == 993) ? 328:
		       /**/
		       (r_counter == 994) ? 329:
		       /**/
		       (r_counter == 995) ? 330:
		       /**/
		       (r_counter == 996) ? 333:
		       /**/
		       (r_counter == 997) ? 334:
		       /**/
		       (r_counter == 998) ? 335:
		       /**/
		       (r_counter == 999) ? 332:
		       /**/
		       (r_counter == 1000) ? 334:
		       /**/
		       (r_counter == 1001) ? 335:
		       /**/
		       (r_counter == 1002) ? 332:
		       /**/
		       (r_counter == 1003) ? 333:
		       /**/
		       (r_counter == 1004) ? 335:
		       /**/
		       (r_counter == 1005) ? 332:
		       /**/
		       (r_counter == 1006) ? 333:
		       /**/
		       (r_counter == 1007) ? 334:
		       /**/
		       (r_counter == 1008) ? 337:
		       /**/
		       (r_counter == 1009) ? 338:
		       /**/
		       (r_counter == 1010) ? 339:
		       /**/
		       (r_counter == 1011) ? 336:
		       /**/
		       (r_counter == 1012) ? 338:
		       /**/
		       (r_counter == 1013) ? 339:
		       /**/
		       (r_counter == 1014) ? 336:
		       /**/
		       (r_counter == 1015) ? 337:
		       /**/
		       (r_counter == 1016) ? 339:
		       /**/
		       (r_counter == 1017) ? 336:
		       /**/
		       (r_counter == 1018) ? 337:
		       /**/
		       (r_counter == 1019) ? 338:
		       /**/
		       (r_counter == 1020) ? 341:
		       /**/
		       (r_counter == 1021) ? 342:
		       /**/
		       (r_counter == 1022) ? 343:
		       /**/
		       (r_counter == 1023) ? 340:
		       /**/
		       (r_counter == 1024) ? 342:
		       /**/
		       (r_counter == 1025) ? 343:
		       /**/
		       (r_counter == 1026) ? 340:
		       /**/
		       (r_counter == 1027) ? 341:
		       /**/
		       (r_counter == 1028) ? 343:
		       /**/
		       (r_counter == 1029) ? 340:
		       /**/
		       (r_counter == 1030) ? 341:
		       /**/
		       (r_counter == 1031) ? 342:
		       /**/
		       (r_counter == 1032) ? 345:
		       /**/
		       (r_counter == 1033) ? 346:
		       /**/
		       (r_counter == 1034) ? 347:
		       /**/
		       (r_counter == 1035) ? 344:
		       /**/
		       (r_counter == 1036) ? 346:
		       /**/
		       (r_counter == 1037) ? 347:
		       /**/
		       (r_counter == 1038) ? 344:
		       /**/
		       (r_counter == 1039) ? 345:
		       /**/
		       (r_counter == 1040) ? 347:
		       /**/
		       (r_counter == 1041) ? 344:
		       /**/
		       (r_counter == 1042) ? 345:
		       /**/
		       (r_counter == 1043) ? 346:
		       /**/
		       (r_counter == 1044) ? 349:
		       /**/
		       (r_counter == 1045) ? 350:
		       /**/
		       (r_counter == 1046) ? 351:
		       /**/
		       (r_counter == 1047) ? 348:
		       /**/
		       (r_counter == 1048) ? 350:
		       /**/
		       (r_counter == 1049) ? 351:
		       /**/
		       (r_counter == 1050) ? 348:
		       /**/
		       (r_counter == 1051) ? 349:
		       /**/
		       (r_counter == 1052) ? 351:
		       /**/
		       (r_counter == 1053) ? 348:
		       /**/
		       (r_counter == 1054) ? 349:
		       /**/
		       (r_counter == 1055) ? 350:
		       /**/
		       (r_counter == 1056) ? 353:
		       /**/
		       (r_counter == 1057) ? 354:
		       /**/
		       (r_counter == 1058) ? 355:
		       /**/
		       (r_counter == 1059) ? 352:
		       /**/
		       (r_counter == 1060) ? 354:
		       /**/
		       (r_counter == 1061) ? 355:
		       /**/
		       (r_counter == 1062) ? 352:
		       /**/
		       (r_counter == 1063) ? 353:
		       /**/
		       (r_counter == 1064) ? 355:
		       /**/
		       (r_counter == 1065) ? 352:
		       /**/
		       (r_counter == 1066) ? 353:
		       /**/
		       (r_counter == 1067) ? 354:
		       /**/
		       (r_counter == 1068) ? 357:
		       /**/
		       (r_counter == 1069) ? 358:
		       /**/
		       (r_counter == 1070) ? 359:
		       /**/
		       (r_counter == 1071) ? 356:
		       /**/
		       (r_counter == 1072) ? 358:
		       /**/
		       (r_counter == 1073) ? 359:
		       /**/
		       (r_counter == 1074) ? 356:
		       /**/
		       (r_counter == 1075) ? 357:
		       /**/
		       (r_counter == 1076) ? 359:
		       /**/
		       (r_counter == 1077) ? 356:
		       /**/
		       (r_counter == 1078) ? 357:
		       /**/
		       (r_counter == 1079) ? 358:
		       /**/
		       (r_counter == 1080) ? 361:
		       /**/
		       (r_counter == 1081) ? 362:
		       /**/
		       (r_counter == 1082) ? 363:
		       /**/
		       (r_counter == 1083) ? 360:
		       /**/
		       (r_counter == 1084) ? 362:
		       /**/
		       (r_counter == 1085) ? 363:
		       /**/
		       (r_counter == 1086) ? 360:
		       /**/
		       (r_counter == 1087) ? 361:
		       /**/
		       (r_counter == 1088) ? 363:
		       /**/
		       (r_counter == 1089) ? 360:
		       /**/
		       (r_counter == 1090) ? 361:
		       /**/
		       (r_counter == 1091) ? 362:
		       /**/
		       (r_counter == 1092) ? 365:
		       /**/
		       (r_counter == 1093) ? 366:
		       /**/
		       (r_counter == 1094) ? 367:
		       /**/
		       (r_counter == 1095) ? 364:
		       /**/
		       (r_counter == 1096) ? 366:
		       /**/
		       (r_counter == 1097) ? 367:
		       /**/
		       (r_counter == 1098) ? 364:
		       /**/
		       (r_counter == 1099) ? 365:
		       /**/
		       (r_counter == 1100) ? 367:
		       /**/
		       (r_counter == 1101) ? 364:
		       /**/
		       (r_counter == 1102) ? 365:
		       /**/
		       (r_counter == 1103) ? 366:
		       /**/
		       (r_counter == 1104) ? 369:
		       /**/
		       (r_counter == 1105) ? 370:
		       /**/
		       (r_counter == 1106) ? 371:
		       /**/
		       (r_counter == 1107) ? 368:
		       /**/
		       (r_counter == 1108) ? 370:
		       /**/
		       (r_counter == 1109) ? 371:
		       /**/
		       (r_counter == 1110) ? 368:
		       /**/
		       (r_counter == 1111) ? 369:
		       /**/
		       (r_counter == 1112) ? 371:
		       /**/
		       (r_counter == 1113) ? 368:
		       /**/
		       (r_counter == 1114) ? 369:
		       /**/
		       (r_counter == 1115) ? 370:
		       /**/
		       (r_counter == 1116) ? 373:
		       /**/
		       (r_counter == 1117) ? 374:
		       /**/
		       (r_counter == 1118) ? 375:
		       /**/
		       (r_counter == 1119) ? 372:
		       /**/
		       (r_counter == 1120) ? 374:
		       /**/
		       (r_counter == 1121) ? 375:
		       /**/
		       (r_counter == 1122) ? 372:
		       /**/
		       (r_counter == 1123) ? 373:
		       /**/
		       (r_counter == 1124) ? 375:
		       /**/
		       (r_counter == 1125) ? 372:
		       /**/
		       (r_counter == 1126) ? 373:
		       /**/
		       (r_counter == 1127) ? 374:
		       /**/
		       (r_counter == 1128) ? 377:
		       /**/
		       (r_counter == 1129) ? 378:
		       /**/
		       (r_counter == 1130) ? 379:
		       /**/
		       (r_counter == 1131) ? 376:
		       /**/
		       (r_counter == 1132) ? 378:
		       /**/
		       (r_counter == 1133) ? 379:
		       /**/
		       (r_counter == 1134) ? 376:
		       /**/
		       (r_counter == 1135) ? 377:
		       /**/
		       (r_counter == 1136) ? 379:
		       /**/
		       (r_counter == 1137) ? 376:
		       /**/
		       (r_counter == 1138) ? 377:
		       /**/
		       (r_counter == 1139) ? 378:
		       /**/
		       (r_counter == 1140) ? 381:
		       /**/
		       (r_counter == 1141) ? 382:
		       /**/
		       (r_counter == 1142) ? 383:
		       /**/
		       (r_counter == 1143) ? 380:
		       /**/
		       (r_counter == 1144) ? 382:
		       /**/
		       (r_counter == 1145) ? 383:
		       /**/
		       (r_counter == 1146) ? 380:
		       /**/
		       (r_counter == 1147) ? 381:
		       /**/
		       (r_counter == 1148) ? 383:
		       /**/
		       (r_counter == 1149) ? 380:
		       /**/
		       (r_counter == 1150) ? 381:
		       /**/
		       (r_counter == 1151) ? 382:
		       /**/
		       (r_counter == 1152) ? 385:
		       /**/
		       (r_counter == 1153) ? 386:
		       /**/
		       (r_counter == 1154) ? 387:
		       /**/
		       (r_counter == 1155) ? 384:
		       /**/
		       (r_counter == 1156) ? 386:
		       /**/
		       (r_counter == 1157) ? 387:
		       /**/
		       (r_counter == 1158) ? 384:
		       /**/
		       (r_counter == 1159) ? 385:
		       /**/
		       (r_counter == 1160) ? 387:
		       /**/
		       (r_counter == 1161) ? 384:
		       /**/
		       (r_counter == 1162) ? 385:
		       /**/
		       (r_counter == 1163) ? 386:
		       /**/
		       (r_counter == 1164) ? 389:
		       /**/
		       (r_counter == 1165) ? 390:
		       /**/
		       (r_counter == 1166) ? 391:
		       /**/
		       (r_counter == 1167) ? 388:
		       /**/
		       (r_counter == 1168) ? 390:
		       /**/
		       (r_counter == 1169) ? 391:
		       /**/
		       (r_counter == 1170) ? 388:
		       /**/
		       (r_counter == 1171) ? 389:
		       /**/
		       (r_counter == 1172) ? 391:
		       /**/
		       (r_counter == 1173) ? 388:
		       /**/
		       (r_counter == 1174) ? 389:
		       /**/
		       (r_counter == 1175) ? 390:
		       /**/
		       (r_counter == 1176) ? 393:
		       /**/
		       (r_counter == 1177) ? 394:
		       /**/
		       (r_counter == 1178) ? 395:
		       /**/
		       (r_counter == 1179) ? 392:
		       /**/
		       (r_counter == 1180) ? 394:
		       /**/
		       (r_counter == 1181) ? 395:
		       /**/
		       (r_counter == 1182) ? 392:
		       /**/
		       (r_counter == 1183) ? 393:
		       /**/
		       (r_counter == 1184) ? 395:
		       /**/
		       (r_counter == 1185) ? 392:
		       /**/
		       (r_counter == 1186) ? 393:
		       /**/
		       (r_counter == 1187) ? 394:
		       /**/
		       (r_counter == 1188) ? 397:
		       /**/
		       (r_counter == 1189) ? 398:
		       /**/
		       (r_counter == 1190) ? 399:
		       /**/
		       (r_counter == 1191) ? 396:
		       /**/
		       (r_counter == 1192) ? 398:
		       /**/
		       (r_counter == 1193) ? 399:
		       /**/
		       (r_counter == 1194) ? 396:
		       /**/
		       (r_counter == 1195) ? 397:
		       /**/
		       (r_counter == 1196) ? 399:
		       /**/
		       (r_counter == 1197) ? 396:
		       /**/
		       (r_counter == 1198) ? 397:
		       /**/
		       (r_counter == 1199) ? 398:
		       /**/
		       (r_counter == 1200) ? 401:
		       /**/
		       (r_counter == 1201) ? 402:
		       /**/
		       (r_counter == 1202) ? 403:
		       /**/
		       (r_counter == 1203) ? 400:
		       /**/
		       (r_counter == 1204) ? 402:
		       /**/
		       (r_counter == 1205) ? 403:
		       /**/
		       (r_counter == 1206) ? 400:
		       /**/
		       (r_counter == 1207) ? 401:
		       /**/
		       (r_counter == 1208) ? 403:
		       /**/
		       (r_counter == 1209) ? 400:
		       /**/
		       (r_counter == 1210) ? 401:
		       /**/
		       (r_counter == 1211) ? 402:
		       /**/
		       (r_counter == 1212) ? 405:
		       /**/
		       (r_counter == 1213) ? 406:
		       /**/
		       (r_counter == 1214) ? 407:
		       /**/
		       (r_counter == 1215) ? 404:
		       /**/
		       (r_counter == 1216) ? 406:
		       /**/
		       (r_counter == 1217) ? 407:
		       /**/
		       (r_counter == 1218) ? 404:
		       /**/
		       (r_counter == 1219) ? 405:
		       /**/
		       (r_counter == 1220) ? 407:
		       /**/
		       (r_counter == 1221) ? 404:
		       /**/
		       (r_counter == 1222) ? 405:
		       /**/
		       (r_counter == 1223) ? 406:
		       /**/
		       (r_counter == 1224) ? 409:
		       /**/
		       (r_counter == 1225) ? 410:
		       /**/
		       (r_counter == 1226) ? 411:
		       /**/
		       (r_counter == 1227) ? 408:
		       /**/
		       (r_counter == 1228) ? 410:
		       /**/
		       (r_counter == 1229) ? 411:
		       /**/
		       (r_counter == 1230) ? 408:
		       /**/
		       (r_counter == 1231) ? 409:
		       /**/
		       (r_counter == 1232) ? 411:
		       /**/
		       (r_counter == 1233) ? 408:
		       /**/
		       (r_counter == 1234) ? 409:
		       /**/
		       (r_counter == 1235) ? 410:
		       /**/
		       (r_counter == 1236) ? 413:
		       /**/
		       (r_counter == 1237) ? 414:
		       /**/
		       (r_counter == 1238) ? 415:
		       /**/
		       (r_counter == 1239) ? 412:
		       /**/
		       (r_counter == 1240) ? 414:
		       /**/
		       (r_counter == 1241) ? 415:
		       /**/
		       (r_counter == 1242) ? 412:
		       /**/
		       (r_counter == 1243) ? 413:
		       /**/
		       (r_counter == 1244) ? 415:
		       /**/
		       (r_counter == 1245) ? 412:
		       /**/
		       (r_counter == 1246) ? 413:
		       /**/
		       (r_counter == 1247) ? 414:
		       /**/
		       (r_counter == 1248) ? 417:
		       /**/
		       (r_counter == 1249) ? 418:
		       /**/
		       (r_counter == 1250) ? 419:
		       /**/
		       (r_counter == 1251) ? 416:
		       /**/
		       (r_counter == 1252) ? 418:
		       /**/
		       (r_counter == 1253) ? 419:
		       /**/
		       (r_counter == 1254) ? 416:
		       /**/
		       (r_counter == 1255) ? 417:
		       /**/
		       (r_counter == 1256) ? 419:
		       /**/
		       (r_counter == 1257) ? 416:
		       /**/
		       (r_counter == 1258) ? 417:
		       /**/
		       (r_counter == 1259) ? 418:
		       /**/
		       (r_counter == 1260) ? 421:
		       /**/
		       (r_counter == 1261) ? 422:
		       /**/
		       (r_counter == 1262) ? 423:
		       /**/
		       (r_counter == 1263) ? 420:
		       /**/
		       (r_counter == 1264) ? 422:
		       /**/
		       (r_counter == 1265) ? 423:
		       /**/
		       (r_counter == 1266) ? 420:
		       /**/
		       (r_counter == 1267) ? 421:
		       /**/
		       (r_counter == 1268) ? 423:
		       /**/
		       (r_counter == 1269) ? 420:
		       /**/
		       (r_counter == 1270) ? 421:
		       /**/
		       (r_counter == 1271) ? 422:
		       /**/
		       (r_counter == 1272) ? 425:
		       /**/
		       (r_counter == 1273) ? 426:
		       /**/
		       (r_counter == 1274) ? 427:
		       /**/
		       (r_counter == 1275) ? 424:
		       /**/
		       (r_counter == 1276) ? 426:
		       /**/
		       (r_counter == 1277) ? 427:
		       /**/
		       (r_counter == 1278) ? 424:
		       /**/
		       (r_counter == 1279) ? 425:
		       /**/
		       (r_counter == 1280) ? 427:
		       /**/
		       (r_counter == 1281) ? 424:
		       /**/
		       (r_counter == 1282) ? 425:
		       /**/
		       (r_counter == 1283) ? 426:
		       /**/
		       (r_counter == 1284) ? 429:
		       /**/
		       (r_counter == 1285) ? 430:
		       /**/
		       (r_counter == 1286) ? 431:
		       /**/
		       (r_counter == 1287) ? 428:
		       /**/
		       (r_counter == 1288) ? 430:
		       /**/
		       (r_counter == 1289) ? 431:
		       /**/
		       (r_counter == 1290) ? 428:
		       /**/
		       (r_counter == 1291) ? 429:
		       /**/
		       (r_counter == 1292) ? 431:
		       /**/
		       (r_counter == 1293) ? 428:
		       /**/
		       (r_counter == 1294) ? 429:
		       /**/
		       (r_counter == 1295) ? 430:
		       /**/
		       (r_counter == 1296) ? 433:
		       /**/
		       (r_counter == 1297) ? 434:
		       /**/
		       (r_counter == 1298) ? 435:
		       /**/
		       (r_counter == 1299) ? 432:
		       /**/
		       (r_counter == 1300) ? 434:
		       /**/
		       (r_counter == 1301) ? 435:
		       /**/
		       (r_counter == 1302) ? 432:
		       /**/
		       (r_counter == 1303) ? 433:
		       /**/
		       (r_counter == 1304) ? 435:
		       /**/
		       (r_counter == 1305) ? 432:
		       /**/
		       (r_counter == 1306) ? 433:
		       /**/
		       (r_counter == 1307) ? 434:
		       /**/
		       (r_counter == 1308) ? 437:
		       /**/
		       (r_counter == 1309) ? 438:
		       /**/
		       (r_counter == 1310) ? 439:
		       /**/
		       (r_counter == 1311) ? 436:
		       /**/
		       (r_counter == 1312) ? 438:
		       /**/
		       (r_counter == 1313) ? 439:
		       /**/
		       (r_counter == 1314) ? 436:
		       /**/
		       (r_counter == 1315) ? 437:
		       /**/
		       (r_counter == 1316) ? 439:
		       /**/
		       (r_counter == 1317) ? 436:
		       /**/
		       (r_counter == 1318) ? 437:
		       /**/
		       (r_counter == 1319) ? 438:
		       /**/
		       (r_counter == 1320) ? 441:
		       /**/
		       (r_counter == 1321) ? 442:
		       /**/
		       (r_counter == 1322) ? 443:
		       /**/
		       (r_counter == 1323) ? 440:
		       /**/
		       (r_counter == 1324) ? 442:
		       /**/
		       (r_counter == 1325) ? 443:
		       /**/
		       (r_counter == 1326) ? 440:
		       /**/
		       (r_counter == 1327) ? 441:
		       /**/
		       (r_counter == 1328) ? 443:
		       /**/
		       (r_counter == 1329) ? 440:
		       /**/
		       (r_counter == 1330) ? 441:
		       /**/
		       (r_counter == 1331) ? 442:
		       /**/
		       (r_counter == 1332) ? 445:
		       /**/
		       (r_counter == 1333) ? 446:
		       /**/
		       (r_counter == 1334) ? 447:
		       /**/
		       (r_counter == 1335) ? 444:
		       /**/
		       (r_counter == 1336) ? 446:
		       /**/
		       (r_counter == 1337) ? 447:
		       /**/
		       (r_counter == 1338) ? 444:
		       /**/
		       (r_counter == 1339) ? 445:
		       /**/
		       (r_counter == 1340) ? 447:
		       /**/
		       (r_counter == 1341) ? 444:
		       /**/
		       (r_counter == 1342) ? 445:
		       /**/
		       (r_counter == 1343) ? 446:
		       /**/
		       (r_counter == 1344) ? 449:
		       /**/
		       (r_counter == 1345) ? 450:
		       /**/
		       (r_counter == 1346) ? 451:
		       /**/
		       (r_counter == 1347) ? 448:
		       /**/
		       (r_counter == 1348) ? 450:
		       /**/
		       (r_counter == 1349) ? 451:
		       /**/
		       (r_counter == 1350) ? 448:
		       /**/
		       (r_counter == 1351) ? 449:
		       /**/
		       (r_counter == 1352) ? 451:
		       /**/
		       (r_counter == 1353) ? 448:
		       /**/
		       (r_counter == 1354) ? 449:
		       /**/
		       (r_counter == 1355) ? 450:
		       /**/
		       (r_counter == 1356) ? 453:
		       /**/
		       (r_counter == 1357) ? 454:
		       /**/
		       (r_counter == 1358) ? 455:
		       /**/
		       (r_counter == 1359) ? 452:
		       /**/
		       (r_counter == 1360) ? 454:
		       /**/
		       (r_counter == 1361) ? 455:
		       /**/
		       (r_counter == 1362) ? 452:
		       /**/
		       (r_counter == 1363) ? 453:
		       /**/
		       (r_counter == 1364) ? 455:
		       /**/
		       (r_counter == 1365) ? 452:
		       /**/
		       (r_counter == 1366) ? 453:
		       /**/
		       (r_counter == 1367) ? 454:
		       /**/
		       (r_counter == 1368) ? 457:
		       /**/
		       (r_counter == 1369) ? 458:
		       /**/
		       (r_counter == 1370) ? 459:
		       /**/
		       (r_counter == 1371) ? 456:
		       /**/
		       (r_counter == 1372) ? 458:
		       /**/
		       (r_counter == 1373) ? 459:
		       /**/
		       (r_counter == 1374) ? 456:
		       /**/
		       (r_counter == 1375) ? 457:
		       /**/
		       (r_counter == 1376) ? 459:
		       /**/
		       (r_counter == 1377) ? 456:
		       /**/
		       (r_counter == 1378) ? 457:
		       /**/
		       (r_counter == 1379) ? 458:
		       /**/
		       (r_counter == 1380) ? 461:
		       /**/
		       (r_counter == 1381) ? 462:
		       /**/
		       (r_counter == 1382) ? 463:
		       /**/
		       (r_counter == 1383) ? 460:
		       /**/
		       (r_counter == 1384) ? 462:
		       /**/
		       (r_counter == 1385) ? 463:
		       /**/
		       (r_counter == 1386) ? 460:
		       /**/
		       (r_counter == 1387) ? 461:
		       /**/
		       (r_counter == 1388) ? 463:
		       /**/
		       (r_counter == 1389) ? 460:
		       /**/
		       (r_counter == 1390) ? 461:
		       /**/
		       (r_counter == 1391) ? 462:
		       /**/
		       (r_counter == 1392) ? 465:
		       /**/
		       (r_counter == 1393) ? 466:
		       /**/
		       (r_counter == 1394) ? 467:
		       /**/
		       (r_counter == 1395) ? 464:
		       /**/
		       (r_counter == 1396) ? 466:
		       /**/
		       (r_counter == 1397) ? 467:
		       /**/
		       (r_counter == 1398) ? 464:
		       /**/
		       (r_counter == 1399) ? 465:
		       /**/
		       (r_counter == 1400) ? 467:
		       /**/
		       (r_counter == 1401) ? 464:
		       /**/
		       (r_counter == 1402) ? 465:
		       /**/
		       (r_counter == 1403) ? 466:
		       /**/
		       (r_counter == 1404) ? 469:
		       /**/
		       (r_counter == 1405) ? 470:
		       /**/
		       (r_counter == 1406) ? 471:
		       /**/
		       (r_counter == 1407) ? 468:
		       /**/
		       (r_counter == 1408) ? 470:
		       /**/
		       (r_counter == 1409) ? 471:
		       /**/
		       (r_counter == 1410) ? 468:
		       /**/
		       (r_counter == 1411) ? 469:
		       /**/
		       (r_counter == 1412) ? 471:
		       /**/
		       (r_counter == 1413) ? 468:
		       /**/
		       (r_counter == 1414) ? 469:
		       /**/
		       (r_counter == 1415) ? 470:
		       /**/
		       (r_counter == 1416) ? 473:
		       /**/
		       (r_counter == 1417) ? 474:
		       /**/
		       (r_counter == 1418) ? 475:
		       /**/
		       (r_counter == 1419) ? 472:
		       /**/
		       (r_counter == 1420) ? 474:
		       /**/
		       (r_counter == 1421) ? 475:
		       /**/
		       (r_counter == 1422) ? 472:
		       /**/
		       (r_counter == 1423) ? 473:
		       /**/
		       (r_counter == 1424) ? 475:
		       /**/
		       (r_counter == 1425) ? 472:
		       /**/
		       (r_counter == 1426) ? 473:
		       /**/
		       (r_counter == 1427) ? 474:
		       /**/
		       (r_counter == 1428) ? 477:
		       /**/
		       (r_counter == 1429) ? 478:
		       /**/
		       (r_counter == 1430) ? 479:
		       /**/
		       (r_counter == 1431) ? 476:
		       /**/
		       (r_counter == 1432) ? 478:
		       /**/
		       (r_counter == 1433) ? 479:
		       /**/
		       (r_counter == 1434) ? 476:
		       /**/
		       (r_counter == 1435) ? 477:
		       /**/
		       (r_counter == 1436) ? 479:
		       /**/
		       (r_counter == 1437) ? 476:
		       /**/
		       (r_counter == 1438) ? 477:
		       /**/
		       (r_counter == 1439) ? 478:
		       /**/
		       (r_counter == 1440) ? 481:
		       /**/
		       (r_counter == 1441) ? 482:
		       /**/
		       (r_counter == 1442) ? 483:
		       /**/
		       (r_counter == 1443) ? 480:
		       /**/
		       (r_counter == 1444) ? 482:
		       /**/
		       (r_counter == 1445) ? 483:
		       /**/
		       (r_counter == 1446) ? 480:
		       /**/
		       (r_counter == 1447) ? 481:
		       /**/
		       (r_counter == 1448) ? 483:
		       /**/
		       (r_counter == 1449) ? 480:
		       /**/
		       (r_counter == 1450) ? 481:
		       /**/
		       (r_counter == 1451) ? 482:
		       /**/
		       (r_counter == 1452) ? 485:
		       /**/
		       (r_counter == 1453) ? 486:
		       /**/
		       (r_counter == 1454) ? 487:
		       /**/
		       (r_counter == 1455) ? 484:
		       /**/
		       (r_counter == 1456) ? 486:
		       /**/
		       (r_counter == 1457) ? 487:
		       /**/
		       (r_counter == 1458) ? 484:
		       /**/
		       (r_counter == 1459) ? 485:
		       /**/
		       (r_counter == 1460) ? 487:
		       /**/
		       (r_counter == 1461) ? 484:
		       /**/
		       (r_counter == 1462) ? 485:
		       /**/
		       (r_counter == 1463) ? 486:
		       /**/
		       (r_counter == 1464) ? 489:
		       /**/
		       (r_counter == 1465) ? 490:
		       /**/
		       (r_counter == 1466) ? 491:
		       /**/
		       (r_counter == 1467) ? 488:
		       /**/
		       (r_counter == 1468) ? 490:
		       /**/
		       (r_counter == 1469) ? 491:
		       /**/
		       (r_counter == 1470) ? 488:
		       /**/
		       (r_counter == 1471) ? 489:
		       /**/
		       (r_counter == 1472) ? 491:
		       /**/
		       (r_counter == 1473) ? 488:
		       /**/
		       (r_counter == 1474) ? 489:
		       /**/
		       (r_counter == 1475) ? 490:
		       /**/
		       (r_counter == 1476) ? 493:
		       /**/
		       (r_counter == 1477) ? 494:
		       /**/
		       (r_counter == 1478) ? 495:
		       /**/
		       (r_counter == 1479) ? 492:
		       /**/
		       (r_counter == 1480) ? 494:
		       /**/
		       (r_counter == 1481) ? 495:
		       /**/
		       (r_counter == 1482) ? 492:
		       /**/
		       (r_counter == 1483) ? 493:
		       /**/
		       (r_counter == 1484) ? 495:
		       /**/
		       (r_counter == 1485) ? 492:
		       /**/
		       (r_counter == 1486) ? 493:
		       /**/
		       (r_counter == 1487) ? 494:
		       /**/
		       (r_counter == 1488) ? 497:
		       /**/
		       (r_counter == 1489) ? 498:
		       /**/
		       (r_counter == 1490) ? 499:
		       /**/
		       (r_counter == 1491) ? 496:
		       /**/
		       (r_counter == 1492) ? 498:
		       /**/
		       (r_counter == 1493) ? 499:
		       /**/
		       (r_counter == 1494) ? 496:
		       /**/
		       (r_counter == 1495) ? 497:
		       /**/
		       (r_counter == 1496) ? 499:
		       /**/
		       (r_counter == 1497) ? 496:
		       /**/
		       (r_counter == 1498) ? 497:
		       /**/
		       (r_counter == 1499) ? 498:
		       /**/
		       (r_counter == 1500) ? 501:
		       /**/
		       (r_counter == 1501) ? 502:
		       /**/
		       (r_counter == 1502) ? 503:
		       /**/
		       (r_counter == 1503) ? 500:
		       /**/
		       (r_counter == 1504) ? 502:
		       /**/
		       (r_counter == 1505) ? 503:
		       /**/
		       (r_counter == 1506) ? 500:
		       /**/
		       (r_counter == 1507) ? 501:
		       /**/
		       (r_counter == 1508) ? 503:
		       /**/
		       (r_counter == 1509) ? 500:
		       /**/
		       (r_counter == 1510) ? 501:
		       /**/
		       (r_counter == 1511) ? 502:
		       /**/
		       (r_counter == 1512) ? 505:
		       /**/
		       (r_counter == 1513) ? 506:
		       /**/
		       (r_counter == 1514) ? 507:
		       /**/
		       (r_counter == 1515) ? 504:
		       /**/
		       (r_counter == 1516) ? 506:
		       /**/
		       (r_counter == 1517) ? 507:
		       /**/
		       (r_counter == 1518) ? 504:
		       /**/
		       (r_counter == 1519) ? 505:
		       /**/
		       (r_counter == 1520) ? 507:
		       /**/
		       (r_counter == 1521) ? 504:
		       /**/
		       (r_counter == 1522) ? 505:
		       /**/
		       (r_counter == 1523) ? 506:
		       /**/
		       (r_counter == 1524) ? 509:
		       /**/
		       (r_counter == 1525) ? 510:
		       /**/
		       (r_counter == 1526) ? 511:
		       /**/
		       (r_counter == 1527) ? 508:
		       /**/
		       (r_counter == 1528) ? 510:
		       /**/
		       (r_counter == 1529) ? 511:
		       /**/
		       (r_counter == 1530) ? 508:
		       /**/
		       (r_counter == 1531) ? 509:
		       /**/
		       (r_counter == 1532) ? 511:
		       /**/
		       (r_counter == 1533) ? 508:
		       /**/
		       (r_counter == 1534) ? 509:
		       /**/
		       (r_counter == 1535) ? 510:
		       /**/
		       (r_counter == 1536) ? 513:
		       /**/
		       (r_counter == 1537) ? 514:
		       /**/
		       (r_counter == 1538) ? 515:
		       /**/
		       (r_counter == 1539) ? 512:
		       /**/
		       (r_counter == 1540) ? 514:
		       /**/
		       (r_counter == 1541) ? 515:
		       /**/
		       (r_counter == 1542) ? 512:
		       /**/
		       (r_counter == 1543) ? 513:
		       /**/
		       (r_counter == 1544) ? 515:
		       /**/
		       (r_counter == 1545) ? 512:
		       /**/
		       (r_counter == 1546) ? 513:
		       /**/
		       (r_counter == 1547) ? 514:
		       /**/
		       (r_counter == 1548) ? 517:
		       /**/
		       (r_counter == 1549) ? 518:
		       /**/
		       (r_counter == 1550) ? 519:
		       /**/
		       (r_counter == 1551) ? 516:
		       /**/
		       (r_counter == 1552) ? 518:
		       /**/
		       (r_counter == 1553) ? 519:
		       /**/
		       (r_counter == 1554) ? 516:
		       /**/
		       (r_counter == 1555) ? 517:
		       /**/
		       (r_counter == 1556) ? 519:
		       /**/
		       (r_counter == 1557) ? 516:
		       /**/
		       (r_counter == 1558) ? 517:
		       /**/
		       (r_counter == 1559) ? 518:
		       /**/
		       (r_counter == 1560) ? 521:
		       /**/
		       (r_counter == 1561) ? 522:
		       /**/
		       (r_counter == 1562) ? 523:
		       /**/
		       (r_counter == 1563) ? 520:
		       /**/
		       (r_counter == 1564) ? 522:
		       /**/
		       (r_counter == 1565) ? 523:
		       /**/
		       (r_counter == 1566) ? 520:
		       /**/
		       (r_counter == 1567) ? 521:
		       /**/
		       (r_counter == 1568) ? 523:
		       /**/
		       (r_counter == 1569) ? 520:
		       /**/
		       (r_counter == 1570) ? 521:
		       /**/
		       (r_counter == 1571) ? 522:
		       /**/
		       (r_counter == 1572) ? 525:
		       /**/
		       (r_counter == 1573) ? 526:
		       /**/
		       (r_counter == 1574) ? 527:
		       /**/
		       (r_counter == 1575) ? 524:
		       /**/
		       (r_counter == 1576) ? 526:
		       /**/
		       (r_counter == 1577) ? 527:
		       /**/
		       (r_counter == 1578) ? 524:
		       /**/
		       (r_counter == 1579) ? 525:
		       /**/
		       (r_counter == 1580) ? 527:
		       /**/
		       (r_counter == 1581) ? 524:
		       /**/
		       (r_counter == 1582) ? 525:
		       /**/
		       (r_counter == 1583) ? 526:
		       /**/
		       (r_counter == 1584) ? 529:
		       /**/
		       (r_counter == 1585) ? 530:
		       /**/
		       (r_counter == 1586) ? 531:
		       /**/
		       (r_counter == 1587) ? 528:
		       /**/
		       (r_counter == 1588) ? 530:
		       /**/
		       (r_counter == 1589) ? 531:
		       /**/
		       (r_counter == 1590) ? 528:
		       /**/
		       (r_counter == 1591) ? 529:
		       /**/
		       (r_counter == 1592) ? 531:
		       /**/
		       (r_counter == 1593) ? 528:
		       /**/
		       (r_counter == 1594) ? 529:
		       /**/
		       (r_counter == 1595) ? 530:
		       /**/
		       (r_counter == 1596) ? 533:
		       /**/
		       (r_counter == 1597) ? 534:
		       /**/
		       (r_counter == 1598) ? 535:
		       /**/
		       (r_counter == 1599) ? 532:
		       /**/
		       (r_counter == 1600) ? 534:
		       /**/
		       (r_counter == 1601) ? 535:
		       /**/
		       (r_counter == 1602) ? 532:
		       /**/
		       (r_counter == 1603) ? 533:
		       /**/
		       (r_counter == 1604) ? 535:
		       /**/
		       (r_counter == 1605) ? 532:
		       /**/
		       (r_counter == 1606) ? 533:
		       /**/
		       (r_counter == 1607) ? 534:
		       /**/
		       (r_counter == 1608) ? 537:
		       /**/
		       (r_counter == 1609) ? 538:
		       /**/
		       (r_counter == 1610) ? 539:
		       /**/
		       (r_counter == 1611) ? 536:
		       /**/
		       (r_counter == 1612) ? 538:
		       /**/
		       (r_counter == 1613) ? 539:
		       /**/
		       (r_counter == 1614) ? 536:
		       /**/
		       (r_counter == 1615) ? 537:
		       /**/
		       (r_counter == 1616) ? 539:
		       /**/
		       (r_counter == 1617) ? 536:
		       /**/
		       (r_counter == 1618) ? 537:
		       /**/
		       (r_counter == 1619) ? 538:
		       /**/
		       (r_counter == 1620) ? 541:
		       /**/
		       (r_counter == 1621) ? 542:
		       /**/
		       (r_counter == 1622) ? 543:
		       /**/
		       (r_counter == 1623) ? 540:
		       /**/
		       (r_counter == 1624) ? 542:
		       /**/
		       (r_counter == 1625) ? 543:
		       /**/
		       (r_counter == 1626) ? 540:
		       /**/
		       (r_counter == 1627) ? 541:
		       /**/
		       (r_counter == 1628) ? 543:
		       /**/
		       (r_counter == 1629) ? 540:
		       /**/
		       (r_counter == 1630) ? 541:
		       /**/
		       (r_counter == 1631) ? 542:
		       /**/
		       (r_counter == 1632) ? 545:
		       /**/
		       (r_counter == 1633) ? 546:
		       /**/
		       (r_counter == 1634) ? 547:
		       /**/
		       (r_counter == 1635) ? 544:
		       /**/
		       (r_counter == 1636) ? 546:
		       /**/
		       (r_counter == 1637) ? 547:
		       /**/
		       (r_counter == 1638) ? 544:
		       /**/
		       (r_counter == 1639) ? 545:
		       /**/
		       (r_counter == 1640) ? 547:
		       /**/
		       (r_counter == 1641) ? 544:
		       /**/
		       (r_counter == 1642) ? 545:
		       /**/
		       (r_counter == 1643) ? 546:
		       /**/
		       (r_counter == 1644) ? 549:
		       /**/
		       (r_counter == 1645) ? 550:
		       /**/
		       (r_counter == 1646) ? 551:
		       /**/
		       (r_counter == 1647) ? 548:
		       /**/
		       (r_counter == 1648) ? 550:
		       /**/
		       (r_counter == 1649) ? 551:
		       /**/
		       (r_counter == 1650) ? 548:
		       /**/
		       (r_counter == 1651) ? 549:
		       /**/
		       (r_counter == 1652) ? 551:
		       /**/
		       (r_counter == 1653) ? 548:
		       /**/
		       (r_counter == 1654) ? 549:
		       /**/
		       (r_counter == 1655) ? 550:
		       /**/
		       (r_counter == 1656) ? 553:
		       /**/
		       (r_counter == 1657) ? 554:
		       /**/
		       (r_counter == 1658) ? 555:
		       /**/
		       (r_counter == 1659) ? 552:
		       /**/
		       (r_counter == 1660) ? 554:
		       /**/
		       (r_counter == 1661) ? 555:
		       /**/
		       (r_counter == 1662) ? 552:
		       /**/
		       (r_counter == 1663) ? 553:
		       /**/
		       (r_counter == 1664) ? 555:
		       /**/
		       (r_counter == 1665) ? 552:
		       /**/
		       (r_counter == 1666) ? 553:
		       /**/
		       (r_counter == 1667) ? 554:
		       /**/
		       (r_counter == 1668) ? 557:
		       /**/
		       (r_counter == 1669) ? 558:
		       /**/
		       (r_counter == 1670) ? 559:
		       /**/
		       (r_counter == 1671) ? 556:
		       /**/
		       (r_counter == 1672) ? 558:
		       /**/
		       (r_counter == 1673) ? 559:
		       /**/
		       (r_counter == 1674) ? 556:
		       /**/
		       (r_counter == 1675) ? 557:
		       /**/
		       (r_counter == 1676) ? 559:
		       /**/
		       (r_counter == 1677) ? 556:
		       /**/
		       (r_counter == 1678) ? 557:
		       /**/
		       (r_counter == 1679) ? 558:
		       /**/
		       (r_counter == 1680) ? 561:
		       /**/
		       (r_counter == 1681) ? 562:
		       /**/
		       (r_counter == 1682) ? 563:
		       /**/
		       (r_counter == 1683) ? 560:
		       /**/
		       (r_counter == 1684) ? 562:
		       /**/
		       (r_counter == 1685) ? 563:
		       /**/
		       (r_counter == 1686) ? 560:
		       /**/
		       (r_counter == 1687) ? 561:
		       /**/
		       (r_counter == 1688) ? 563:
		       /**/
		       (r_counter == 1689) ? 560:
		       /**/
		       (r_counter == 1690) ? 561:
		       /**/
		       (r_counter == 1691) ? 562:
		       /**/
		       (r_counter == 1692) ? 565:
		       /**/
		       (r_counter == 1693) ? 566:
		       /**/
		       (r_counter == 1694) ? 567:
		       /**/
		       (r_counter == 1695) ? 564:
		       /**/
		       (r_counter == 1696) ? 566:
		       /**/
		       (r_counter == 1697) ? 567:
		       /**/
		       (r_counter == 1698) ? 564:
		       /**/
		       (r_counter == 1699) ? 565:
		       /**/
		       (r_counter == 1700) ? 567:
		       /**/
		       (r_counter == 1701) ? 564:
		       /**/
		       (r_counter == 1702) ? 565:
		       /**/
		       (r_counter == 1703) ? 566:
		       /**/
		       (r_counter == 1704) ? 569:
		       /**/
		       (r_counter == 1705) ? 570:
		       /**/
		       (r_counter == 1706) ? 571:
		       /**/
		       (r_counter == 1707) ? 568:
		       /**/
		       (r_counter == 1708) ? 570:
		       /**/
		       (r_counter == 1709) ? 571:
		       /**/
		       (r_counter == 1710) ? 568:
		       /**/
		       (r_counter == 1711) ? 569:
		       /**/
		       (r_counter == 1712) ? 571:
		       /**/
		       (r_counter == 1713) ? 568:
		       /**/
		       (r_counter == 1714) ? 569:
		       /**/
		       (r_counter == 1715) ? 570:
		       /**/
		       (r_counter == 1716) ? 573:
		       /**/
		       (r_counter == 1717) ? 574:
		       /**/
		       (r_counter == 1718) ? 575:
		       /**/
		       (r_counter == 1719) ? 572:
		       /**/
		       (r_counter == 1720) ? 574:
		       /**/
		       (r_counter == 1721) ? 575:
		       /**/
		       (r_counter == 1722) ? 572:
		       /**/
		       (r_counter == 1723) ? 573:
		       /**/
		       (r_counter == 1724) ? 575:
		       /**/
		       (r_counter == 1725) ? 572:
		       /**/
		       (r_counter == 1726) ? 573:
		       /**/
		       (r_counter == 1727) ? 574:
		       /**/
		       (r_counter == 1728) ? 577:
		       /**/
		       (r_counter == 1729) ? 578:
		       /**/
		       (r_counter == 1730) ? 579:
		       /**/
		       (r_counter == 1731) ? 576:
		       /**/
		       (r_counter == 1732) ? 578:
		       /**/
		       (r_counter == 1733) ? 579:
		       /**/
		       (r_counter == 1734) ? 576:
		       /**/
		       (r_counter == 1735) ? 577:
		       /**/
		       (r_counter == 1736) ? 579:
		       /**/
		       (r_counter == 1737) ? 576:
		       /**/
		       (r_counter == 1738) ? 577:
		       /**/
		       (r_counter == 1739) ? 578:
		       /**/
		       (r_counter == 1740) ? 581:
		       /**/
		       (r_counter == 1741) ? 582:
		       /**/
		       (r_counter == 1742) ? 583:
		       /**/
		       (r_counter == 1743) ? 580:
		       /**/
		       (r_counter == 1744) ? 582:
		       /**/
		       (r_counter == 1745) ? 583:
		       /**/
		       (r_counter == 1746) ? 580:
		       /**/
		       (r_counter == 1747) ? 581:
		       /**/
		       (r_counter == 1748) ? 583:
		       /**/
		       (r_counter == 1749) ? 580:
		       /**/
		       (r_counter == 1750) ? 581:
		       /**/
		       (r_counter == 1751) ? 582:
		       /**/
		       (r_counter == 1752) ? 585:
		       /**/
		       (r_counter == 1753) ? 586:
		       /**/
		       (r_counter == 1754) ? 587:
		       /**/
		       (r_counter == 1755) ? 584:
		       /**/
		       (r_counter == 1756) ? 586:
		       /**/
		       (r_counter == 1757) ? 587:
		       /**/
		       (r_counter == 1758) ? 584:
		       /**/
		       (r_counter == 1759) ? 585:
		       /**/
		       (r_counter == 1760) ? 587:
		       /**/
		       (r_counter == 1761) ? 584:
		       /**/
		       (r_counter == 1762) ? 585:
		       /**/
		       (r_counter == 1763) ? 586:
		       /**/
		       (r_counter == 1764) ? 589:
		       /**/
		       (r_counter == 1765) ? 590:
		       /**/
		       (r_counter == 1766) ? 591:
		       /**/
		       (r_counter == 1767) ? 588:
		       /**/
		       (r_counter == 1768) ? 590:
		       /**/
		       (r_counter == 1769) ? 591:
		       /**/
		       (r_counter == 1770) ? 588:
		       /**/
		       (r_counter == 1771) ? 589:
		       /**/
		       (r_counter == 1772) ? 591:
		       /**/
		       (r_counter == 1773) ? 588:
		       /**/
		       (r_counter == 1774) ? 589:
		       /**/
		       (r_counter == 1775) ? 590:
		       /**/
		       (r_counter == 1776) ? 593:
		       /**/
		       (r_counter == 1777) ? 594:
		       /**/
		       (r_counter == 1778) ? 595:
		       /**/
		       (r_counter == 1779) ? 592:
		       /**/
		       (r_counter == 1780) ? 594:
		       /**/
		       (r_counter == 1781) ? 595:
		       /**/
		       (r_counter == 1782) ? 592:
		       /**/
		       (r_counter == 1783) ? 593:
		       /**/
		       (r_counter == 1784) ? 595:
		       /**/
		       (r_counter == 1785) ? 592:
		       /**/
		       (r_counter == 1786) ? 593:
		       /**/
		       (r_counter == 1787) ? 594:
		       /**/
		       (r_counter == 1788) ? 597:
		       /**/
		       (r_counter == 1789) ? 598:
		       /**/
		       (r_counter == 1790) ? 599:
		       /**/
		       (r_counter == 1791) ? 596:
		       /**/
		       (r_counter == 1792) ? 598:
		       /**/
		       (r_counter == 1793) ? 599:
		       /**/
		       (r_counter == 1794) ? 596:
		       /**/
		       (r_counter == 1795) ? 597:
		       /**/
		       (r_counter == 1796) ? 599:
		       /**/
		       (r_counter == 1797) ? 596:
		       /**/
		       (r_counter == 1798) ? 597:
		       /**/
		       (r_counter == 1799) ? 598:
		       /**/
		       (r_counter == 1800) ? 601:
		       /**/
		       (r_counter == 1801) ? 602:
		       /**/
		       (r_counter == 1802) ? 603:
		       /**/
		       (r_counter == 1803) ? 600:
		       /**/
		       (r_counter == 1804) ? 602:
		       /**/
		       (r_counter == 1805) ? 603:
		       /**/
		       (r_counter == 1806) ? 600:
		       /**/
		       (r_counter == 1807) ? 601:
		       /**/
		       (r_counter == 1808) ? 603:
		       /**/
		       (r_counter == 1809) ? 600:
		       /**/
		       (r_counter == 1810) ? 601:
		       /**/
		       (r_counter == 1811) ? 602:
		       /**/
		       (r_counter == 1812) ? 605:
		       /**/
		       (r_counter == 1813) ? 606:
		       /**/
		       (r_counter == 1814) ? 607:
		       /**/
		       (r_counter == 1815) ? 604:
		       /**/
		       (r_counter == 1816) ? 606:
		       /**/
		       (r_counter == 1817) ? 607:
		       /**/
		       (r_counter == 1818) ? 604:
		       /**/
		       (r_counter == 1819) ? 605:
		       /**/
		       (r_counter == 1820) ? 607:
		       /**/
		       (r_counter == 1821) ? 604:
		       /**/
		       (r_counter == 1822) ? 605:
		       /**/
		       (r_counter == 1823) ? 606:
		       /**/
		       (r_counter == 1824) ? 609:
		       /**/
		       (r_counter == 1825) ? 610:
		       /**/
		       (r_counter == 1826) ? 611:
		       /**/
		       (r_counter == 1827) ? 608:
		       /**/
		       (r_counter == 1828) ? 610:
		       /**/
		       (r_counter == 1829) ? 611:
		       /**/
		       (r_counter == 1830) ? 608:
		       /**/
		       (r_counter == 1831) ? 609:
		       /**/
		       (r_counter == 1832) ? 611:
		       /**/
		       (r_counter == 1833) ? 608:
		       /**/
		       (r_counter == 1834) ? 609:
		       /**/
		       (r_counter == 1835) ? 610:
		       /**/
		       (r_counter == 1836) ? 613:
		       /**/
		       (r_counter == 1837) ? 614:
		       /**/
		       (r_counter == 1838) ? 615:
		       /**/
		       (r_counter == 1839) ? 612:
		       /**/
		       (r_counter == 1840) ? 614:
		       /**/
		       (r_counter == 1841) ? 615:
		       /**/
		       (r_counter == 1842) ? 612:
		       /**/
		       (r_counter == 1843) ? 613:
		       /**/
		       (r_counter == 1844) ? 615:
		       /**/
		       (r_counter == 1845) ? 612:
		       /**/
		       (r_counter == 1846) ? 613:
		       /**/
		       (r_counter == 1847) ? 614:
		       /**/
		       (r_counter == 1848) ? 617:
		       /**/
		       (r_counter == 1849) ? 618:
		       /**/
		       (r_counter == 1850) ? 619:
		       /**/
		       (r_counter == 1851) ? 616:
		       /**/
		       (r_counter == 1852) ? 618:
		       /**/
		       (r_counter == 1853) ? 619:
		       /**/
		       (r_counter == 1854) ? 616:
		       /**/
		       (r_counter == 1855) ? 617:
		       /**/
		       (r_counter == 1856) ? 619:
		       /**/
		       (r_counter == 1857) ? 616:
		       /**/
		       (r_counter == 1858) ? 617:
		       /**/
		       (r_counter == 1859) ? 618:
		       /**/
		       (r_counter == 1860) ? 621:
		       /**/
		       (r_counter == 1861) ? 622:
		       /**/
		       (r_counter == 1862) ? 623:
		       /**/
		       (r_counter == 1863) ? 620:
		       /**/
		       (r_counter == 1864) ? 622:
		       /**/
		       (r_counter == 1865) ? 623:
		       /**/
		       (r_counter == 1866) ? 620:
		       /**/
		       (r_counter == 1867) ? 621:
		       /**/
		       (r_counter == 1868) ? 623:
		       /**/
		       (r_counter == 1869) ? 620:
		       /**/
		       (r_counter == 1870) ? 621:
		       /**/
		       (r_counter == 1871) ? 622:
		       /**/
		       (r_counter == 1872) ? 625:
		       /**/
		       (r_counter == 1873) ? 626:
		       /**/
		       (r_counter == 1874) ? 627:
		       /**/
		       (r_counter == 1875) ? 624:
		       /**/
		       (r_counter == 1876) ? 626:
		       /**/
		       (r_counter == 1877) ? 627:
		       /**/
		       (r_counter == 1878) ? 624:
		       /**/
		       (r_counter == 1879) ? 625:
		       /**/
		       (r_counter == 1880) ? 627:
		       /**/
		       (r_counter == 1881) ? 624:
		       /**/
		       (r_counter == 1882) ? 625:
		       /**/
		       (r_counter == 1883) ? 626:
		       /**/
		       (r_counter == 1884) ? 629:
		       /**/
		       (r_counter == 1885) ? 630:
		       /**/
		       (r_counter == 1886) ? 631:
		       /**/
		       (r_counter == 1887) ? 628:
		       /**/
		       (r_counter == 1888) ? 630:
		       /**/
		       (r_counter == 1889) ? 631:
		       /**/
		       (r_counter == 1890) ? 628:
		       /**/
		       (r_counter == 1891) ? 629:
		       /**/
		       (r_counter == 1892) ? 631:
		       /**/
		       (r_counter == 1893) ? 628:
		       /**/
		       (r_counter == 1894) ? 629:
		       /**/
		       (r_counter == 1895) ? 630:
		       /**/
		       (r_counter == 1896) ? 633:
		       /**/
		       (r_counter == 1897) ? 634:
		       /**/
		       (r_counter == 1898) ? 635:
		       /**/
		       (r_counter == 1899) ? 632:
		       /**/
		       (r_counter == 1900) ? 634:
		       /**/
		       (r_counter == 1901) ? 635:
		       /**/
		       (r_counter == 1902) ? 632:
		       /**/
		       (r_counter == 1903) ? 633:
		       /**/
		       (r_counter == 1904) ? 635:
		       /**/
		       (r_counter == 1905) ? 632:
		       /**/
		       (r_counter == 1906) ? 633:
		       /**/
		       (r_counter == 1907) ? 634:
		       /**/
		       (r_counter == 1908) ? 637:
		       /**/
		       (r_counter == 1909) ? 638:
		       /**/
		       (r_counter == 1910) ? 639:
		       /**/
		       (r_counter == 1911) ? 636:
		       /**/
		       (r_counter == 1912) ? 638:
		       /**/
		       (r_counter == 1913) ? 639:
		       /**/
		       (r_counter == 1914) ? 636:
		       /**/
		       (r_counter == 1915) ? 637:
		       /**/
		       (r_counter == 1916) ? 639:
		       /**/
		       (r_counter == 1917) ? 636:
		       /**/
		       (r_counter == 1918) ? 637:
		       /**/
		       (r_counter == 1919) ? 638:
		       /**/
		       (r_counter == 1920) ? 641:
		       /**/
		       (r_counter == 1921) ? 642:
		       /**/
		       (r_counter == 1922) ? 643:
		       /**/
		       (r_counter == 1923) ? 640:
		       /**/
		       (r_counter == 1924) ? 642:
		       /**/
		       (r_counter == 1925) ? 643:
		       /**/
		       (r_counter == 1926) ? 640:
		       /**/
		       (r_counter == 1927) ? 641:
		       /**/
		       (r_counter == 1928) ? 643:
		       /**/
		       (r_counter == 1929) ? 640:
		       /**/
		       (r_counter == 1930) ? 641:
		       /**/
		       (r_counter == 1931) ? 642:
		       /**/
		       (r_counter == 1932) ? 645:
		       /**/
		       (r_counter == 1933) ? 646:
		       /**/
		       (r_counter == 1934) ? 647:
		       /**/
		       (r_counter == 1935) ? 644:
		       /**/
		       (r_counter == 1936) ? 646:
		       /**/
		       (r_counter == 1937) ? 647:
		       /**/
		       (r_counter == 1938) ? 644:
		       /**/
		       (r_counter == 1939) ? 645:
		       /**/
		       (r_counter == 1940) ? 647:
		       /**/
		       (r_counter == 1941) ? 644:
		       /**/
		       (r_counter == 1942) ? 645:
		       /**/
		       (r_counter == 1943) ? 646:
		       /**/
		       (r_counter == 1944) ? 649:
		       /**/
		       (r_counter == 1945) ? 650:
		       /**/
		       (r_counter == 1946) ? 651:
		       /**/
		       (r_counter == 1947) ? 648:
		       /**/
		       (r_counter == 1948) ? 650:
		       /**/
		       (r_counter == 1949) ? 651:
		       /**/
		       (r_counter == 1950) ? 648:
		       /**/
		       (r_counter == 1951) ? 649:
		       /**/
		       (r_counter == 1952) ? 651:
		       /**/
		       (r_counter == 1953) ? 648:
		       /**/
		       (r_counter == 1954) ? 649:
		       /**/
		       (r_counter == 1955) ? 650:
		       /**/
		       (r_counter == 1956) ? 653:
		       /**/
		       (r_counter == 1957) ? 654:
		       /**/
		       (r_counter == 1958) ? 655:
		       /**/
		       (r_counter == 1959) ? 652:
		       /**/
		       (r_counter == 1960) ? 654:
		       /**/
		       (r_counter == 1961) ? 655:
		       /**/
		       (r_counter == 1962) ? 652:
		       /**/
		       (r_counter == 1963) ? 653:
		       /**/
		       (r_counter == 1964) ? 655:
		       /**/
		       (r_counter == 1965) ? 652:
		       /**/
		       (r_counter == 1966) ? 653:
		       /**/
		       (r_counter == 1967) ? 654:
		       /**/
		       (r_counter == 1968) ? 657:
		       /**/
		       (r_counter == 1969) ? 658:
		       /**/
		       (r_counter == 1970) ? 659:
		       /**/
		       (r_counter == 1971) ? 656:
		       /**/
		       (r_counter == 1972) ? 658:
		       /**/
		       (r_counter == 1973) ? 659:
		       /**/
		       (r_counter == 1974) ? 656:
		       /**/
		       (r_counter == 1975) ? 657:
		       /**/
		       (r_counter == 1976) ? 659:
		       /**/
		       (r_counter == 1977) ? 656:
		       /**/
		       (r_counter == 1978) ? 657:
		       /**/
		       (r_counter == 1979) ? 658:
		       /**/
		       (r_counter == 1980) ? 661:
		       /**/
		       (r_counter == 1981) ? 662:
		       /**/
		       (r_counter == 1982) ? 663:
		       /**/
		       (r_counter == 1983) ? 660:
		       /**/
		       (r_counter == 1984) ? 662:
		       /**/
		       (r_counter == 1985) ? 663:
		       /**/
		       (r_counter == 1986) ? 660:
		       /**/
		       (r_counter == 1987) ? 661:
		       /**/
		       (r_counter == 1988) ? 663:
		       /**/
		       (r_counter == 1989) ? 660:
		       /**/
		       (r_counter == 1990) ? 661:
		       /**/
		       (r_counter == 1991) ? 662:
		       /**/
		       (r_counter == 1992) ? 665:
		       /**/
		       (r_counter == 1993) ? 666:
		       /**/
		       (r_counter == 1994) ? 667:
		       /**/
		       (r_counter == 1995) ? 664:
		       /**/
		       (r_counter == 1996) ? 666:
		       /**/
		       (r_counter == 1997) ? 667:
		       /**/
		       (r_counter == 1998) ? 664:
		       /**/
		       (r_counter == 1999) ? 665:
		       /**/
		       (r_counter == 2000) ? 667:
		       /**/
		       (r_counter == 2001) ? 664:
		       /**/
		       (r_counter == 2002) ? 665:
		       /**/
		       (r_counter == 2003) ? 666:
		       /**/
		       (r_counter == 2004) ? 669:
		       /**/
		       (r_counter == 2005) ? 670:
		       /**/
		       (r_counter == 2006) ? 671:
		       /**/
		       (r_counter == 2007) ? 668:
		       /**/
		       (r_counter == 2008) ? 670:
		       /**/
		       (r_counter == 2009) ? 671:
		       /**/
		       (r_counter == 2010) ? 668:
		       /**/
		       (r_counter == 2011) ? 669:
		       /**/
		       (r_counter == 2012) ? 671:
		       /**/
		       (r_counter == 2013) ? 668:
		       /**/
		       (r_counter == 2014) ? 669:
		       /**/
		       (r_counter == 2015) ? 670:
		       /**/
		       (r_counter == 2016) ? 673:
		       /**/
		       (r_counter == 2017) ? 674:
		       /**/
		       (r_counter == 2018) ? 675:
		       /**/
		       (r_counter == 2019) ? 672:
		       /**/
		       (r_counter == 2020) ? 674:
		       /**/
		       (r_counter == 2021) ? 675:
		       /**/
		       (r_counter == 2022) ? 672:
		       /**/
		       (r_counter == 2023) ? 673:
		       /**/
		       (r_counter == 2024) ? 675:
		       /**/
		       (r_counter == 2025) ? 672:
		       /**/
		       (r_counter == 2026) ? 673:
		       /**/
		       (r_counter == 2027) ? 674:
		       /**/
		       (r_counter == 2028) ? 677:
		       /**/
		       (r_counter == 2029) ? 678:
		       /**/
		       (r_counter == 2030) ? 679:
		       /**/
		       (r_counter == 2031) ? 676:
		       /**/
		       (r_counter == 2032) ? 678:
		       /**/
		       (r_counter == 2033) ? 679:
		       /**/
		       (r_counter == 2034) ? 676:
		       /**/
		       (r_counter == 2035) ? 677:
		       /**/
		       (r_counter == 2036) ? 679:
		       /**/
		       (r_counter == 2037) ? 676:
		       /**/
		       (r_counter == 2038) ? 677:
		       /**/
		       (r_counter == 2039) ? 678:
		       /**/
		       (r_counter == 2040) ? 681:
		       /**/
		       (r_counter == 2041) ? 682:
		       /**/
		       (r_counter == 2042) ? 683:
		       /**/
		       (r_counter == 2043) ? 680:
		       /**/
		       (r_counter == 2044) ? 682:
		       /**/
		       (r_counter == 2045) ? 683:
		       /**/
		       (r_counter == 2046) ? 680:
		       /**/
		       (r_counter == 2047) ? 681:
		       /**/
		       (r_counter == 2048) ? 683:
		       /**/
		       (r_counter == 2049) ? 680:
		       /**/
		       (r_counter == 2050) ? 681:
		       /**/
		       (r_counter == 2051) ? 682:
		       /**/
		       (r_counter == 2052) ? 685:
		       /**/
		       (r_counter == 2053) ? 686:
		       /**/
		       (r_counter == 2054) ? 687:
		       /**/
		       (r_counter == 2055) ? 684:
		       /**/
		       (r_counter == 2056) ? 686:
		       /**/
		       (r_counter == 2057) ? 687:
		       /**/
		       (r_counter == 2058) ? 684:
		       /**/
		       (r_counter == 2059) ? 685:
		       /**/
		       (r_counter == 2060) ? 687:
		       /**/
		       (r_counter == 2061) ? 684:
		       /**/
		       (r_counter == 2062) ? 685:
		       /**/
		       (r_counter == 2063) ? 686:
		       /**/
		       (r_counter == 2064) ? 689:
		       /**/
		       (r_counter == 2065) ? 690:
		       /**/
		       (r_counter == 2066) ? 691:
		       /**/
		       (r_counter == 2067) ? 688:
		       /**/
		       (r_counter == 2068) ? 690:
		       /**/
		       (r_counter == 2069) ? 691:
		       /**/
		       (r_counter == 2070) ? 688:
		       /**/
		       (r_counter == 2071) ? 689:
		       /**/
		       (r_counter == 2072) ? 691:
		       /**/
		       (r_counter == 2073) ? 688:
		       /**/
		       (r_counter == 2074) ? 689:
		       /**/
		       (r_counter == 2075) ? 690:
		       /**/
		       (r_counter == 2076) ? 693:
		       /**/
		       (r_counter == 2077) ? 694:
		       /**/
		       (r_counter == 2078) ? 695:
		       /**/
		       (r_counter == 2079) ? 692:
		       /**/
		       (r_counter == 2080) ? 694:
		       /**/
		       (r_counter == 2081) ? 695:
		       /**/
		       (r_counter == 2082) ? 692:
		       /**/
		       (r_counter == 2083) ? 693:
		       /**/
		       (r_counter == 2084) ? 695:
		       /**/
		       (r_counter == 2085) ? 692:
		       /**/
		       (r_counter == 2086) ? 693:
		       /**/
		       (r_counter == 2087) ? 694:
		       /**/
		       (r_counter == 2088) ? 697:
		       /**/
		       (r_counter == 2089) ? 698:
		       /**/
		       (r_counter == 2090) ? 699:
		       /**/
		       (r_counter == 2091) ? 696:
		       /**/
		       (r_counter == 2092) ? 698:
		       /**/
		       (r_counter == 2093) ? 699:
		       /**/
		       (r_counter == 2094) ? 696:
		       /**/
		       (r_counter == 2095) ? 697:
		       /**/
		       (r_counter == 2096) ? 699:
		       /**/
		       (r_counter == 2097) ? 696:
		       /**/
		       (r_counter == 2098) ? 697:
		       /**/
		       (r_counter == 2099) ? 698:
		       /**/
		       (r_counter == 2100) ? 701:
		       /**/
		       (r_counter == 2101) ? 702:
		       /**/
		       (r_counter == 2102) ? 703:
		       /**/
		       (r_counter == 2103) ? 700:
		       /**/
		       (r_counter == 2104) ? 702:
		       /**/
		       (r_counter == 2105) ? 703:
		       /**/
		       (r_counter == 2106) ? 700:
		       /**/
		       (r_counter == 2107) ? 701:
		       /**/
		       (r_counter == 2108) ? 703:
		       /**/
		       (r_counter == 2109) ? 700:
		       /**/
		       (r_counter == 2110) ? 701:
		       /**/
		       (r_counter == 2111) ? 702:
		       /**/
		       (r_counter == 2112) ? 705:
		       /**/
		       (r_counter == 2113) ? 706:
		       /**/
		       (r_counter == 2114) ? 707:
		       /**/
		       (r_counter == 2115) ? 704:
		       /**/
		       (r_counter == 2116) ? 706:
		       /**/
		       (r_counter == 2117) ? 707:
		       /**/
		       (r_counter == 2118) ? 704:
		       /**/
		       (r_counter == 2119) ? 705:
		       /**/
		       (r_counter == 2120) ? 707:
		       /**/
		       (r_counter == 2121) ? 704:
		       /**/
		       (r_counter == 2122) ? 705:
		       /**/
		       (r_counter == 2123) ? 706:
		       /**/
		       (r_counter == 2124) ? 709:
		       /**/
		       (r_counter == 2125) ? 710:
		       /**/
		       (r_counter == 2126) ? 711:
		       /**/
		       (r_counter == 2127) ? 708:
		       /**/
		       (r_counter == 2128) ? 710:
		       /**/
		       (r_counter == 2129) ? 711:
		       /**/
		       (r_counter == 2130) ? 708:
		       /**/
		       (r_counter == 2131) ? 709:
		       /**/
		       (r_counter == 2132) ? 711:
		       /**/
		       (r_counter == 2133) ? 708:
		       /**/
		       (r_counter == 2134) ? 709:
		       /**/
		       (r_counter == 2135) ? 710:
		       /**/
		       (r_counter == 2136) ? 713:
		       /**/
		       (r_counter == 2137) ? 714:
		       /**/
		       (r_counter == 2138) ? 715:
		       /**/
		       (r_counter == 2139) ? 712:
		       /**/
		       (r_counter == 2140) ? 714:
		       /**/
		       (r_counter == 2141) ? 715:
		       /**/
		       (r_counter == 2142) ? 712:
		       /**/
		       (r_counter == 2143) ? 713:
		       /**/
		       (r_counter == 2144) ? 715:
		       /**/
		       (r_counter == 2145) ? 712:
		       /**/
		       (r_counter == 2146) ? 713:
		       /**/
		       (r_counter == 2147) ? 714:
		       /**/
		       (r_counter == 2148) ? 717:
		       /**/
		       (r_counter == 2149) ? 718:
		       /**/
		       (r_counter == 2150) ? 719:
		       /**/
		       (r_counter == 2151) ? 716:
		       /**/
		       (r_counter == 2152) ? 718:
		       /**/
		       (r_counter == 2153) ? 719:
		       /**/
		       (r_counter == 2154) ? 716:
		       /**/
		       (r_counter == 2155) ? 717:
		       /**/
		       (r_counter == 2156) ? 719:
		       /**/
		       (r_counter == 2157) ? 716:
		       /**/
		       (r_counter == 2158) ? 717:
		       /**/
		       (r_counter == 2159) ? 718:
		       /**/
		       (r_counter == 2160) ? 721:
		       /**/
		       (r_counter == 2161) ? 722:
		       /**/
		       (r_counter == 2162) ? 723:
		       /**/
		       (r_counter == 2163) ? 720:
		       /**/
		       (r_counter == 2164) ? 722:
		       /**/
		       (r_counter == 2165) ? 723:
		       /**/
		       (r_counter == 2166) ? 720:
		       /**/
		       (r_counter == 2167) ? 721:
		       /**/
		       (r_counter == 2168) ? 723:
		       /**/
		       (r_counter == 2169) ? 720:
		       /**/
		       (r_counter == 2170) ? 721:
		       /**/
		       (r_counter == 2171) ? 722:
		       /**/
		       (r_counter == 2172) ? 725:
		       /**/
		       (r_counter == 2173) ? 726:
		       /**/
		       (r_counter == 2174) ? 727:
		       /**/
		       (r_counter == 2175) ? 724:
		       /**/
		       (r_counter == 2176) ? 726:
		       /**/
		       (r_counter == 2177) ? 727:
		       /**/
		       (r_counter == 2178) ? 724:
		       /**/
		       (r_counter == 2179) ? 725:
		       /**/
		       (r_counter == 2180) ? 727:
		       /**/
		       (r_counter == 2181) ? 724:
		       /**/
		       (r_counter == 2182) ? 725:
		       /**/
		       (r_counter == 2183) ? 726:
		       /**/
		       (r_counter == 2184) ? 729:
		       /**/
		       (r_counter == 2185) ? 730:
		       /**/
		       (r_counter == 2186) ? 731:
		       /**/
		       (r_counter == 2187) ? 728:
		       /**/
		       (r_counter == 2188) ? 730:
		       /**/
		       (r_counter == 2189) ? 731:
		       /**/
		       (r_counter == 2190) ? 728:
		       /**/
		       (r_counter == 2191) ? 729:
		       /**/
		       (r_counter == 2192) ? 731:
		       /**/
		       (r_counter == 2193) ? 728:
		       /**/
		       (r_counter == 2194) ? 729:
		       /**/
		       (r_counter == 2195) ? 730:
		       /**/
		       (r_counter == 2196) ? 733:
		       /**/
		       (r_counter == 2197) ? 734:
		       /**/
		       (r_counter == 2198) ? 735:
		       /**/
		       (r_counter == 2199) ? 732:
		       /**/
		       (r_counter == 2200) ? 734:
		       /**/
		       (r_counter == 2201) ? 735:
		       /**/
		       (r_counter == 2202) ? 732:
		       /**/
		       (r_counter == 2203) ? 733:
		       /**/
		       (r_counter == 2204) ? 735:
		       /**/
		       (r_counter == 2205) ? 732:
		       /**/
		       (r_counter == 2206) ? 733:
		       /**/
		       (r_counter == 2207) ? 734:
		       /**/
		       (r_counter == 2208) ? 737:
		       /**/
		       (r_counter == 2209) ? 738:
		       /**/
		       (r_counter == 2210) ? 739:
		       /**/
		       (r_counter == 2211) ? 736:
		       /**/
		       (r_counter == 2212) ? 738:
		       /**/
		       (r_counter == 2213) ? 739:
		       /**/
		       (r_counter == 2214) ? 736:
		       /**/
		       (r_counter == 2215) ? 737:
		       /**/
		       (r_counter == 2216) ? 739:
		       /**/
		       (r_counter == 2217) ? 736:
		       /**/
		       (r_counter == 2218) ? 737:
		       /**/
		       (r_counter == 2219) ? 738:
		       /**/
		       (r_counter == 2220) ? 741:
		       /**/
		       (r_counter == 2221) ? 742:
		       /**/
		       (r_counter == 2222) ? 743:
		       /**/
		       (r_counter == 2223) ? 740:
		       /**/
		       (r_counter == 2224) ? 742:
		       /**/
		       (r_counter == 2225) ? 743:
		       /**/
		       (r_counter == 2226) ? 740:
		       /**/
		       (r_counter == 2227) ? 741:
		       /**/
		       (r_counter == 2228) ? 743:
		       /**/
		       (r_counter == 2229) ? 740:
		       /**/
		       (r_counter == 2230) ? 741:
		       /**/
		       (r_counter == 2231) ? 742:
		       /**/
		       (r_counter == 2232) ? 745:
		       /**/
		       (r_counter == 2233) ? 746:
		       /**/
		       (r_counter == 2234) ? 747:
		       /**/
		       (r_counter == 2235) ? 744:
		       /**/
		       (r_counter == 2236) ? 746:
		       /**/
		       (r_counter == 2237) ? 747:
		       /**/
		       (r_counter == 2238) ? 744:
		       /**/
		       (r_counter == 2239) ? 745:
		       /**/
		       (r_counter == 2240) ? 747:
		       /**/
		       (r_counter == 2241) ? 744:
		       /**/
		       (r_counter == 2242) ? 745:
		       /**/
		       (r_counter == 2243) ? 746:
		       /**/
		       (r_counter == 2244) ? 749:
		       /**/
		       (r_counter == 2245) ? 750:
		       /**/
		       (r_counter == 2246) ? 751:
		       /**/
		       (r_counter == 2247) ? 748:
		       /**/
		       (r_counter == 2248) ? 750:
		       /**/
		       (r_counter == 2249) ? 751:
		       /**/
		       (r_counter == 2250) ? 748:
		       /**/
		       (r_counter == 2251) ? 749:
		       /**/
		       (r_counter == 2252) ? 751:
		       /**/
		       (r_counter == 2253) ? 748:
		       /**/
		       (r_counter == 2254) ? 749:
		       /**/
		       (r_counter == 2255) ? 750:
		       /**/
		       (r_counter == 2256) ? 753:
		       /**/
		       (r_counter == 2257) ? 754:
		       /**/
		       (r_counter == 2258) ? 755:
		       /**/
		       (r_counter == 2259) ? 752:
		       /**/
		       (r_counter == 2260) ? 754:
		       /**/
		       (r_counter == 2261) ? 755:
		       /**/
		       (r_counter == 2262) ? 752:
		       /**/
		       (r_counter == 2263) ? 753:
		       /**/
		       (r_counter == 2264) ? 755:
		       /**/
		       (r_counter == 2265) ? 752:
		       /**/
		       (r_counter == 2266) ? 753:
		       /**/
		       (r_counter == 2267) ? 754:
		       /**/
		       (r_counter == 2268) ? 757:
		       /**/
		       (r_counter == 2269) ? 758:
		       /**/
		       (r_counter == 2270) ? 759:
		       /**/
		       (r_counter == 2271) ? 756:
		       /**/
		       (r_counter == 2272) ? 758:
		       /**/
		       (r_counter == 2273) ? 759:
		       /**/
		       (r_counter == 2274) ? 756:
		       /**/
		       (r_counter == 2275) ? 757:
		       /**/
		       (r_counter == 2276) ? 759:
		       /**/
		       (r_counter == 2277) ? 756:
		       /**/
		       (r_counter == 2278) ? 757:
		       /**/
		       (r_counter == 2279) ? 758:
		       /**/
		       (r_counter == 2280) ? 761:
		       /**/
		       (r_counter == 2281) ? 762:
		       /**/
		       (r_counter == 2282) ? 763:
		       /**/
		       (r_counter == 2283) ? 760:
		       /**/
		       (r_counter == 2284) ? 762:
		       /**/
		       (r_counter == 2285) ? 763:
		       /**/
		       (r_counter == 2286) ? 760:
		       /**/
		       (r_counter == 2287) ? 761:
		       /**/
		       (r_counter == 2288) ? 763:
		       /**/
		       (r_counter == 2289) ? 760:
		       /**/
		       (r_counter == 2290) ? 761:
		       /**/
		       (r_counter == 2291) ? 762:
		       /**/
		       (r_counter == 2292) ? 765:
		       /**/
		       (r_counter == 2293) ? 766:
		       /**/
		       (r_counter == 2294) ? 767:
		       /**/
		       (r_counter == 2295) ? 764:
		       /**/
		       (r_counter == 2296) ? 766:
		       /**/
		       (r_counter == 2297) ? 767:
		       /**/
		       (r_counter == 2298) ? 764:
		       /**/
		       (r_counter == 2299) ? 765:
		       /**/
		       (r_counter == 2300) ? 767:
		       /**/
		       (r_counter == 2301) ? 764:
		       /**/
		       (r_counter == 2302) ? 765:
		       /**/
		       (r_counter == 2303) ? 766:
		       /**/
		       (r_counter == 2304) ? 769:
		       /**/
		       (r_counter == 2305) ? 770:
		       /**/
		       (r_counter == 2306) ? 771:
		       /**/
		       (r_counter == 2307) ? 768:
		       /**/
		       (r_counter == 2308) ? 770:
		       /**/
		       (r_counter == 2309) ? 771:
		       /**/
		       (r_counter == 2310) ? 768:
		       /**/
		       (r_counter == 2311) ? 769:
		       /**/
		       (r_counter == 2312) ? 771:
		       /**/
		       (r_counter == 2313) ? 768:
		       /**/
		       (r_counter == 2314) ? 769:
		       /**/
		       (r_counter == 2315) ? 770:
		       /**/
		       (r_counter == 2316) ? 773:
		       /**/
		       (r_counter == 2317) ? 774:
		       /**/
		       (r_counter == 2318) ? 775:
		       /**/
		       (r_counter == 2319) ? 772:
		       /**/
		       (r_counter == 2320) ? 774:
		       /**/
		       (r_counter == 2321) ? 775:
		       /**/
		       (r_counter == 2322) ? 772:
		       /**/
		       (r_counter == 2323) ? 773:
		       /**/
		       (r_counter == 2324) ? 775:
		       /**/
		       (r_counter == 2325) ? 772:
		       /**/
		       (r_counter == 2326) ? 773:
		       /**/
		       (r_counter == 2327) ? 774:
		       /**/
		       (r_counter == 2328) ? 777:
		       /**/
		       (r_counter == 2329) ? 778:
		       /**/
		       (r_counter == 2330) ? 779:
		       /**/
		       (r_counter == 2331) ? 776:
		       /**/
		       (r_counter == 2332) ? 778:
		       /**/
		       (r_counter == 2333) ? 779:
		       /**/
		       (r_counter == 2334) ? 776:
		       /**/
		       (r_counter == 2335) ? 777:
		       /**/
		       (r_counter == 2336) ? 779:
		       /**/
		       (r_counter == 2337) ? 776:
		       /**/
		       (r_counter == 2338) ? 777:
		       /**/
		       (r_counter == 2339) ? 778:
		       /**/
		       (r_counter == 2340) ? 781:
		       /**/
		       (r_counter == 2341) ? 782:
		       /**/
		       (r_counter == 2342) ? 783:
		       /**/
		       (r_counter == 2343) ? 780:
		       /**/
		       (r_counter == 2344) ? 782:
		       /**/
		       (r_counter == 2345) ? 783:
		       /**/
		       (r_counter == 2346) ? 780:
		       /**/
		       (r_counter == 2347) ? 781:
		       /**/
		       (r_counter == 2348) ? 783:
		       /**/
		       (r_counter == 2349) ? 780:
		       /**/
		       (r_counter == 2350) ? 781:
		       /**/
		       (r_counter == 2351) ? 782:
		       /**/
		       (r_counter == 2352) ? 785:
		       /**/
		       (r_counter == 2353) ? 786:
		       /**/
		       (r_counter == 2354) ? 787:
		       /**/
		       (r_counter == 2355) ? 784:
		       /**/
		       (r_counter == 2356) ? 786:
		       /**/
		       (r_counter == 2357) ? 787:
		       /**/
		       (r_counter == 2358) ? 784:
		       /**/
		       (r_counter == 2359) ? 785:
		       /**/
		       (r_counter == 2360) ? 787:
		       /**/
		       (r_counter == 2361) ? 784:
		       /**/
		       (r_counter == 2362) ? 785:
		       /**/
		       (r_counter == 2363) ? 786:
		       /**/
		       (r_counter == 2364) ? 789:
		       /**/
		       (r_counter == 2365) ? 790:
		       /**/
		       (r_counter == 2366) ? 791:
		       /**/
		       (r_counter == 2367) ? 788:
		       /**/
		       (r_counter == 2368) ? 790:
		       /**/
		       (r_counter == 2369) ? 791:
		       /**/
		       (r_counter == 2370) ? 788:
		       /**/
		       (r_counter == 2371) ? 789:
		       /**/
		       (r_counter == 2372) ? 791:
		       /**/
		       (r_counter == 2373) ? 788:
		       /**/
		       (r_counter == 2374) ? 789:
		       /**/
		       (r_counter == 2375) ? 790:
		       /**/
		       (r_counter == 2376) ? 793:
		       /**/
		       (r_counter == 2377) ? 794:
		       /**/
		       (r_counter == 2378) ? 795:
		       /**/
		       (r_counter == 2379) ? 792:
		       /**/
		       (r_counter == 2380) ? 794:
		       /**/
		       (r_counter == 2381) ? 795:
		       /**/
		       (r_counter == 2382) ? 792:
		       /**/
		       (r_counter == 2383) ? 793:
		       /**/
		       (r_counter == 2384) ? 795:
		       /**/
		       (r_counter == 2385) ? 792:
		       /**/
		       (r_counter == 2386) ? 793:
		       /**/
		       (r_counter == 2387) ? 794:
		       /**/
		       (r_counter == 2388) ? 797:
		       /**/
		       (r_counter == 2389) ? 798:
		       /**/
		       (r_counter == 2390) ? 799:
		       /**/
		       (r_counter == 2391) ? 796:
		       /**/
		       (r_counter == 2392) ? 798:
		       /**/
		       (r_counter == 2393) ? 799:
		       /**/
		       (r_counter == 2394) ? 796:
		       /**/
		       (r_counter == 2395) ? 797:
		       /**/
		       (r_counter == 2396) ? 799:
		       /**/
		       (r_counter == 2397) ? 796:
		       /**/
		       (r_counter == 2398) ? 797:
		       /**/
		       (r_counter == 2399) ? 798:
		       /**/
		       0;
   assign i_wdata_beta=(r_state == zStateBetaInit) ? o_rdata_lambda:
		       (r_state == zStateColumn) ? o_data_test_beta:
		       0;

   assign o_column_data = 
			  /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 2) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 3 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 4) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 5 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 6) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 7 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 8) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 9 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 10) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 11 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 12) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 13 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 14) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 15 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 16) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 17 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 18) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 19 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 20) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 21 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 22) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 23 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 24) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 25 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 26) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 27 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 28) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 29 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 30) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 31 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 32) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 33 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 34) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 35 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 36) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 37 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 38) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 39 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 40) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 41 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 42) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 43 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 44) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 45 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 46) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 47 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 48) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 49 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 50) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 51 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 52) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 53 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 54) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 55 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 56) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 57 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 58) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 59 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 60) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 61 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 62) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 63 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 64) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 65 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 66) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 67 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 68) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 69 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 70) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 71 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 72) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 73 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 74) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 75 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 76) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 77 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 78) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 79 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 80) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 81 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 82) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 83 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 84) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 85 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 86) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 87 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 88) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 89 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 90) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 91 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 92) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 93 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 94) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 95 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 96) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 97 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 98) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 99 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 100) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 101 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 102) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 103 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 104) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 105 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 106) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 107 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 108) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 109 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 110) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 111 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 112) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 113 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 114) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 115 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 116) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 117 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 118) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 119 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 120) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 121 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 122) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 123 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 124) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 125 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 126) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 127 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 128) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 129 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 130) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 131 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 132) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 133 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 134) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 135 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 136) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 137 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 138) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 139 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 140) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 141 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 142) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 143 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 144) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 145 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 146) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 147 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 148) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 149 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 150) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 151 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 152) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 153 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 154) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 155 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 156) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 157 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 158) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 159 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 160) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 161 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 162) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 163 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 164) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 165 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 166) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 167 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 168) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 169 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 170) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 171 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 172) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 173 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 174) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 175 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 176) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 177 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 178) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 179 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 180) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 181 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 182) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 183 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 184) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 185 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 186) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 187 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 188) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 189 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 190) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 191 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 192) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 193 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 194) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 195 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 196) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 197 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 198) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 199 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 200) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 201 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 202) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 203 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 204) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 205 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 206) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 207 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 208) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 209 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 210) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 211 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 212) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 213 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 214) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 215 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 216) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 217 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 218) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 219 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 220) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 221 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 222) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 223 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 224) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 225 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 226) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 227 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 228) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 229 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 230) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 231 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 232) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 233 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 234) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 235 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 236) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 237 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 238) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 239 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 240) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 241 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 242) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 243 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 244) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 245 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 246) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 247 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 248) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 249 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 250) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 251 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 252) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 253 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 254) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 255 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 256) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 257 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 258) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 259 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 260) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 261 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 262) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 263 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 264) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 265 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 266) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 267 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 268) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 269 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 270) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 271 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 272) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 273 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 274) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 275 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 276) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 277 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 278) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 279 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 280) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 281 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 282) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 283 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 284) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 285 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 286) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 287 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 288) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 289 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 290) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 291 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 292) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 293 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 294) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 295 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 296) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 297 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 298) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 299 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 300) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 301 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 302) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 303 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 304) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 305 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 306) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 307 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 308) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 309 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 310) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 311 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 312) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 313 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 314) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 315 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 316) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 317 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 318) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 319 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 320) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 321 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 322) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 323 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 324) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 325 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 326) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 327 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 328) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 329 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 330) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 331 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 332) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 333 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 334) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 335 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 336) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 337 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 338) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 339 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 340) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 341 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 342) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 343 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 344) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 345 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 346) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 347 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 348) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 349 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 350) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 351 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 352) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 353 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 354) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 355 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 356) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 357 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 358) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 359 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 360) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 361 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 362) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 363 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 364) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 365 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 366) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 367 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 368) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 369 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 370) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 371 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 372) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 373 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 374) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 375 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 376) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 377 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 378) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 379 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 380) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 381 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 382) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 383 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 384) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 385 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 386) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 387 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 388) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 389 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 390) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 391 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 392) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 393 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 394) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 395 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 396) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 397 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 398) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 399 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 400) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 401 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 402) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 403 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 404) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 405 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 406) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 407 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 408) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 409 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 410) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 411 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 412) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 413 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 414) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 415 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 416) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 417 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 418) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 419 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 420) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 421 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 422) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 423 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 424) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 425 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 426) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 427 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 428) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 429 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 430) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 431 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 432) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 433 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 434) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 435 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 436) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 437 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 438) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 439 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 440) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 441 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 442) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 443 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 444) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 445 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 446) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 447 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 448) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 449 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 450) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 451 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 452) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 453 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 454) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 455 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 456) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 457 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 458) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 459 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 460) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 461 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 462) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 463 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 464) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 465 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 466) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 467 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 468) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 469 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 470) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 471 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 472) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 473 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 474) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 475 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 476) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 477 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 478) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 479 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 480) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 481 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 482) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 483 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 484) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 485 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 486) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 487 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 488) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 489 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 490) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 491 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 492) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 493 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 494) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 495 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 496) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 497 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 498) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 499 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 500) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 501 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 502) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 503 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 504) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 505 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 506) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 507 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 508) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 509 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 510) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 511 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 512) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 513 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 514) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 515 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 516) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 517 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 518) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 519 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 520) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 521 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 522) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 523 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 524) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 525 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 526) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 527 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 528) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 529 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 530) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 531 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 532) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 533 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 534) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 535 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 536) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 537 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 538) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 539 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 540) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 541 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 542) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 543 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 544) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 545 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 546) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 547 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 548) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 549 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 550) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 551 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 552) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 553 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 554) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 555 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 556) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 557 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 558) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 559 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 560) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 561 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 562) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 563 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 564) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 565 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 566) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 567 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 568) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 569 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 570) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 571 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 572) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 573 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 574) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 575 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 576) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 577 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 578) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 579 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 580) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 581 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 582) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 583 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 584) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 585 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 586) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 587 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 588) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 589 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 590) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 591 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 592) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 593 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 594) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 595 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 596) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 597 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 598) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 599 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 600) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 601 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 602) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 603 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 604) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 605 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 606) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 607 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 608) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 609 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 610) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 611 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 612) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 613 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 614) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 615 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 616) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 617 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 618) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 619 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 620) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 621 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 622) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 623 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 624) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 625 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 626) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 627 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 628) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 629 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 630) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 631 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 632) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 633 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 634) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 635 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 636) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 637 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 638) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 639 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 640) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 641 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 642) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 643 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 644) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 645 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 646) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 647 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 648) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 649 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 650) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 651 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 652) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 653 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 654) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 655 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 656) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 657 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 658) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 659 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 660) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 661 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 662) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 663 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 664) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 665 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 666) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 667 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 668) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 669 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 670) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 671 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 672) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 673 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 674) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 675 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 676) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 677 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 678) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 679 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 680) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 681 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 682) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 683 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 684) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 685 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 686) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 687 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 688) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 689 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 690) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 691 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 692) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 693 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 694) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 695 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 696) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 697 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 698) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 699 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 700) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 701 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 702) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 703 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 704) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 705 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 706) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 707 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 708) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 709 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 710) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 711 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 712) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 713 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 714) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 715 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 716) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 717 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 718) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 719 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 720) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 721 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 722) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 723 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 724) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 725 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 726) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 727 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 728) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 729 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 730) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 731 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 732) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 733 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 734) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 735 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 736) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 737 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 738) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 739 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 740) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 741 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 742) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 743 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 744) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 745 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 746) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 747 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 748) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 749 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 750) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 751 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 752) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 753 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 754) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 755 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 756) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 757 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 758) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 759 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 760) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 761 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 762) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 763 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 764) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 765 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 766) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 767 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 768) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 769 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 770) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 771 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 772) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 773 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 774) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 775 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 776) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 777 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 778) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 779 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 780) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 781 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 782) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 783 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 784) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 785 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 786) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 787 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 788) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 789 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 790) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 791 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 792) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 793 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 794) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 795 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 796) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 797 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 798) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 799 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 800) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 801 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 802) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 803 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 804) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 805 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 806) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 807 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 808) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 809 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 810) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 811 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 812) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 813 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 814) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 815 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 816) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 817 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 818) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 819 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 820) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 821 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 822) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 823 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 824) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 825 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 826) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 827 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 828) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 829 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 830) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 831 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 832) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 833 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 834) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 835 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 836) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 837 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 838) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 839 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 840) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 841 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 842) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 843 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 844) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 845 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 846) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 847 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 848) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 849 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 850) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 851 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 852) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 853 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 854) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 855 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 856) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 857 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 858) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 859 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 860) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 861 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 862) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 863 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 864) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 865 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 866) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 867 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 868) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 869 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 870) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 871 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 872) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 873 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 874) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 875 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 876) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 877 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 878) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 879 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 880) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 881 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 882) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 883 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 884) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 885 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 886) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 887 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 888) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 889 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 890) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 891 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 892) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 893 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 894) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 895 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 896) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 897 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 898) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 899 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 900) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 901 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 902) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 903 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 904) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 905 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 906) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 907 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 908) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 909 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 910) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 911 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 912) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 913 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 914) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 915 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 916) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 917 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 918) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 919 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 920) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 921 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 922) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 923 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 924) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 925 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 926) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 927 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 928) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 929 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 930) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 931 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 932) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 933 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 934) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 935 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 936) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 937 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 938) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 939 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 940) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 941 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 942) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 943 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 944) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 945 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 946) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 947 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 948) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 949 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 950) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 951 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 952) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 953 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 954) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 955 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 956) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 957 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 958) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 959 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 960) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 961 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 962) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 963 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 964) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 965 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 966) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 967 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 968) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 969 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 970) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 971 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 972) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 973 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 974) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 975 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 976) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 977 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 978) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 979 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 980) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 981 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 982) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 983 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 984) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 985 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 986) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 987 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 988) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 989 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 990) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 991 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 992) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 993 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 994) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 995 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 996) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 997 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 998) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 999 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1000) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1001 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1002) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1003 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1004) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1005 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1006) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1007 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1008) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1009 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1010) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1011 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1012) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1013 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1014) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1015 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1016) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1017 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1018) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1019 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1020) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1021 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1022) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1023 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1024) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1025 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1026) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1027 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1028) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1029 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1030) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1031 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1032) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1033 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1034) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1035 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1036) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1037 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1038) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1039 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1040) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1041 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1042) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1043 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1044) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1045 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1046) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1047 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1048) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1049 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1050) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1051 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1052) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1053 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1054) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1055 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1056) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1057 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1058) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1059 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1060) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1061 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1062) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1063 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1064) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1065 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1066) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1067 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1068) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1069 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1070) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1071 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1072) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1073 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1074) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1075 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1076) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1077 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1078) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1079 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1080) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1081 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1082) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1083 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1084) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1085 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1086) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1087 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1088) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1089 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1090) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1091 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1092) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1093 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1094) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1095 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1096) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1097 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1098) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1099 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1100) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1101 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1102) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1103 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1104) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1105 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1106) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1107 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1108) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1109 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1110) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1111 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1112) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1113 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1114) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1115 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1116) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1117 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1118) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1119 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1120) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1121 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1122) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1123 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1124) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1125 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1126) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1127 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1128) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1129 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1130) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1131 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1132) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1133 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1134) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1135 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1136) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1137 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1138) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1139 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1140) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1141 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1142) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1143 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1144) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1145 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1146) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1147 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1148) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1149 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1150) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1151 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1152) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1153 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1154) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1155 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1156) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1157 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1158) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1159 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1160) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1161 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1162) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1163 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1164) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1165 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1166) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1167 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1168) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1169 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1170) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1171 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1172) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1173 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1174) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1175 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1176) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1177 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1178) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1179 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1180) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1181 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1182) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1183 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1184) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1185 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1186) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1187 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1188) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1189 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1190) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1191 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1192) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1193 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1194) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1195 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1196) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1197 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1198) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1199 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1200) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1201 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1202) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1203 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1204) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1205 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1206) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1207 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1208) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1209 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1210) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1211 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1212) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1213 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1214) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1215 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1216) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1217 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1218) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1219 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1220) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1221 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1222) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1223 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1224) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1225 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1226) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1227 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1228) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1229 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1230) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1231 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1232) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1233 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1234) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1235 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1236) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1237 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1238) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1239 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1240) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1241 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1242) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1243 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1244) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1245 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1246) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1247 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1248) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1249 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1250) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1251 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1252) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1253 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1254) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1255 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1256) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1257 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1258) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1259 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1260) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1261 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1262) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1263 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1264) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1265 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1266) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1267 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1268) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1269 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1270) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1271 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1272) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1273 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1274) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1275 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1276) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1277 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1278) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1279 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1280) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1281 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1282) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1283 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1284) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1285 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1286) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1287 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1288) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1289 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1290) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1291 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1292) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1293 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1294) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1295 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1296) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1297 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1298) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1299 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1300) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1301 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1302) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1303 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1304) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1305 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1306) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1307 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1308) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1309 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1310) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1311 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1312) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1313 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1314) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1315 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1316) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1317 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1318) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1319 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1320) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1321 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1322) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1323 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1324) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1325 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1326) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1327 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1328) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1329 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1330) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1331 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1332) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1333 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1334) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1335 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1336) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1337 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1338) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1339 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1340) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1341 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1342) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1343 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1344) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1345 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1346) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1347 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1348) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1349 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1350) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1351 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1352) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1353 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1354) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1355 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1356) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1357 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1358) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1359 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1360) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1361 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1362) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1363 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1364) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1365 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1366) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1367 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1368) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1369 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1370) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1371 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1372) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1373 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1374) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1375 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1376) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1377 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1378) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1379 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1380) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1381 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1382) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1383 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1384) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1385 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1386) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1387 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1388) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1389 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1390) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1391 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1392) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1393 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1394) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1395 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1396) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1397 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1398) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1399 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1400) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1401 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1402) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1403 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1404) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1405 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1406) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1407 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1408) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1409 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1410) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1411 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1412) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1413 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1414) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1415 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1416) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1417 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1418) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1419 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1420) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1421 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1422) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1423 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1424) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1425 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1426) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1427 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1428) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1429 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1430) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1431 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1432) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1433 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1434) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1435 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1436) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1437 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1438) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1439 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1440) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1441 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1442) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1443 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1444) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1445 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1446) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1447 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1448) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1449 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1450) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1451 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1452) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1453 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1454) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1455 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1456) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1457 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1458) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1459 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1460) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1461 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1462) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1463 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1464) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1465 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1466) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1467 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1468) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1469 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1470) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1471 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1472) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1473 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1474) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1475 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1476) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1477 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1478) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1479 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1480) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1481 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1482) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1483 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1484) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1485 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1486) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1487 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1488) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1489 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1490) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1491 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1492) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1493 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1494) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1495 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1496) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1497 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1498) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1499 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1500) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1501 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1502) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1503 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1504) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1505 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1506) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1507 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1508) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1509 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1510) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1511 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1512) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1513 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1514) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1515 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1516) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1517 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1518) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1519 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1520) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1521 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1522) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1523 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1524) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1525 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1526) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1527 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1528) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1529 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1530) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1531 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1532) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1533 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1534) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1535 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1536) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1537 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1538) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1539 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1540) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1541 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1542) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1543 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1544) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1545 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1546) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1547 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1548) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1549 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1550) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1551 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1552) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1553 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1554) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1555 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1556) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1557 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1558) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1559 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1560) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1561 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1562) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1563 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1564) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1565 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1566) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1567 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1568) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1569 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1570) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1571 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1572) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1573 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1574) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1575 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1576) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1577 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1578) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1579 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1580) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1581 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1582) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1583 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1584) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1585 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1586) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1587 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1588) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1589 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1590) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1591 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1592) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1593 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1594) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1595 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1596) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1597 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1598) ? o_rdata_lambda:
			  /**/
				    /**/
			  /**/
			  (r_state == zStateColumn) &(r_counter == 1599 ) ? o_rdata_alpha:
				    /**/
				    /**/
			  /**/ 
			  (r_state == zStateColumn) & (r_counter == 1600) ? o_rdata_lambda:
			  /**/
				    /**/
				    /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 2 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 3) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 4 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 5 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 6) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 7 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 8 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 9) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 10 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 11 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 12) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 13 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 14 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 15) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 16 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 17 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 18) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 19 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 20 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 21) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 22 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 23 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 24) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 25 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 26 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 27) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 28 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 29 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 30) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 31 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 32 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 33) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 34 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 35 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 36) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 37 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 38 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 39) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 40 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 41 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 42) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 43 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 44 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 45) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 46 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 47 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 48) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 49 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 50 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 51) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 52 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 53 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 54) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 55 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 56 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 57) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 58 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 59 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 60) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 61 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 62 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 63) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 64 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 65 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 66) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 67 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 68 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 69) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 70 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 71 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 72) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 73 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 74 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 75) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 76 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 77 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 78) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 79 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 80 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 81) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 82 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 83 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 84) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 85 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 86 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 87) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 88 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 89 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 90) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 91 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 92 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 93) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 94 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 95 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 96) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 97 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 98 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 99) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 100 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 101 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 102) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 103 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 104 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 105) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 106 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 107 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 108) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 109 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 110 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 111) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 112 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 113 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 114) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 115 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 116 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 117) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 118 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 119 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 120) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 121 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 122 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 123) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 124 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 125 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 126) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 127 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 128 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 129) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 130 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 131 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 132) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 133 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 134 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 135) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 136 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 137 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 138) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 139 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 140 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 141) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 142 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 143 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 144) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 145 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 146 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 147) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 148 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 149 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 150) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 151 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 152 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 153) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 154 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 155 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 156) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 157 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 158 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 159) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 160 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 161 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 162) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 163 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 164 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 165) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 166 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 167 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 168) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 169 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 170 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 171) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 172 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 173 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 174) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 175 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 176 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 177) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 178 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 179 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 180) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 181 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 182 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 183) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 184 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 185 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 186) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 187 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 188 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 189) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 190 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 191 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 192) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 193 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 194 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 195) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 196 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 197 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 198) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 199 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 200 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 201) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 202 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 203 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 204) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 205 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 206 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 207) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 208 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 209 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 210) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 211 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 212 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 213) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 214 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 215 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 216) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 217 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 218 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 219) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 220 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 221 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 222) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 223 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 224 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 225) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 226 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 227 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 228) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 229 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 230 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 231) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 232 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 233 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 234) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 235 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 236 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 237) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 238 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 239 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 240) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 241 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 242 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 243) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 244 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 245 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 246) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 247 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 248 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 249) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 250 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 251 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 252) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 253 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 254 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 255) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 256 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 257 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 258) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 259 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 260 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 261) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 262 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 263 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 264) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 265 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 266 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 267) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 268 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 269 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 270) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 271 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 272 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 273) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 274 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 275 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 276) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 277 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 278 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 279) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 280 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 281 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 282) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 283 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 284 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 285) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 286 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 287 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 288) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 289 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 290 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 291) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 292 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 293 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 294) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 295 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 296 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 297) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 298 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 299 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 300) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 301 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 302 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 303) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 304 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 305 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 306) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 307 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 308 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 309) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 310 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 311 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 312) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 313 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 314 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 315) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 316 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 317 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 318) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 319 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 320 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 321) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 322 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 323 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 324) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 325 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 326 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 327) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 328 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 329 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 330) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 331 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 332 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 333) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 334 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 335 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 336) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 337 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 338 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 339) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 340 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 341 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 342) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 343 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 344 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 345) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 346 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 347 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 348) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 349 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 350 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 351) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 352 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 353 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 354) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 355 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 356 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 357) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 358 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 359 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 360) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 361 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 362 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 363) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 364 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 365 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 366) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 367 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 368 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 369) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 370 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 371 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 372) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 373 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 374 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 375) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 376 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 377 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 378) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 379 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 380 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 381) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 382 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 383 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 384) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 385 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 386 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 387) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 388 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 389 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 390) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 391 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 392 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 393) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 394 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 395 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 396) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 397 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 398 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 399) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 400 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 401 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 402) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 403 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 404 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 405) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 406 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 407 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 408) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 409 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 410 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 411) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 412 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 413 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 414) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 415 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 416 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 417) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 418 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 419 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 420) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 421 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 422 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 423) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 424 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 425 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 426) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 427 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 428 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 429) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 430 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 431 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 432) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 433 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 434 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 435) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 436 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 437 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 438) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 439 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 440 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 441) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 442 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 443 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 444) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 445 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 446 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 447) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 448 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 449 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 450) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 451 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 452 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 453) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 454 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 455 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 456) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 457 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 458 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 459) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 460 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 461 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 462) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 463 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 464 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 465) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 466 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 467 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 468) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 469 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 470 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 471) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 472 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 473 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 474) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 475 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 476 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 477) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 478 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 479 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 480) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 481 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 482 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 483) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 484 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 485 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 486) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 487 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 488 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 489) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 490 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 491 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 492) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 493 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 494 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 495) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 496 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 497 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 498) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 499 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 500 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 501) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 502 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 503 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 504) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 505 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 506 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 507) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 508 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 509 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 510) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 511 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 512 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 513) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 514 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 515 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 516) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 517 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 518 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 519) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 520 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 521 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 522) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 523 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 524 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 525) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 526 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 527 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 528) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 529 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 530 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 531) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 532 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 533 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 534) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 535 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 536 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 537) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 538 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 539 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 540) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 541 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 542 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 543) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 544 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 545 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 546) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 547 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 548 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 549) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 550 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 551 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 552) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 553 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 554 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 555) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 556 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 557 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 558) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 559 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 560 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 561) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 562 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 563 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 564) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 565 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 566 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 567) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 568 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 569 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 570) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 571 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 572 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 573) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 574 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 575 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 576) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 577 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 578 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 579) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 580 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 581 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 582) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 583 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 584 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 585) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 586 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 587 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 588) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 589 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 590 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 591) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 592 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 593 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 594) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 595 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 596 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 597) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 598 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 599 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 600) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 601 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 602 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 603) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 604 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 605 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 606) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 607 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 608 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 609) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 610 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 611 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 612) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 613 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 614 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 615) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 616 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 617 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 618) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 619 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 620 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 621) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 622 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 623 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 624) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 625 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 626 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 627) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 628 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 629 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 630) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 631 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 632 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 633) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 634 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 635 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 636) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 637 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 638 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 639) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 640 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 641 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 642) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 643 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 644 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 645) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 646 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 647 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 648) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 649 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 650 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 651) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 652 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 653 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 654) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 655 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 656 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 657) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 658 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 659 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 660) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 661 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 662 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 663) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 664 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 665 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 666) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 667 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 668 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 669) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 670 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 671 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 672) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 673 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 674 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 675) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 676 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 677 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 678) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 679 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 680 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 681) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 682 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 683 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 684) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 685 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 686 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 687) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 688 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 689 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 690) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 691 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 692 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 693) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 694 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 695 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 696) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 697 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 698 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 699) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 700 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 701 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 702) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 703 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 704 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 705) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 706 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 707 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 708) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 709 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 710 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 711) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 712 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 713 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 714) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 715 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 716 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 717) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 718 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 719 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 720) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 721 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 722 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 723) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 724 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 725 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 726) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 727 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 728 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 729) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 730 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 731 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 732) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 733 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 734 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 735) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 736 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 737 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 738) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 739 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 740 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 741) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 742 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 743 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 744) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 745 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 746 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 747) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 748 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 749 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 750) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 751 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 752 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 753) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 754 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 755 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 756) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 757 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 758 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 759) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 760 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 761 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 762) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 763 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 764 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 765) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 766 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 767 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 768) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 769 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 770 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 771) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 772 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 773 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 774) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 775 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 776 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 777) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 778 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 779 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 780) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 781 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 782 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 783) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 784 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 785 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 786) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 787 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 788 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 789) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 790 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 791 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 792) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 793 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 794 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 795) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 796 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 797 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 798) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 799 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 800 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 801) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 802 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 803 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 804) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 805 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 806 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 807) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 808 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 809 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 810) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 811 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 812 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 813) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 814 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 815 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 816) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 817 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 818 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 819) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 820 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 821 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 822) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 823 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 824 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 825) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 826 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 827 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 828) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 829 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 830 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 831) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 832 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 833 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 834) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 835 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 836 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 837) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 838 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 839 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 840) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 841 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 842 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 843) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 844 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 845 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 846) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 847 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 848 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 849) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 850 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 851 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 852) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 853 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 854 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 855) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 856 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 857 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 858) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 859 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 860 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 861) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 862 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 863 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 864) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 865 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 866 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 867) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 868 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 869 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 870) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 871 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 872 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 873) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 874 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 875 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 876) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 877 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 878 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 879) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 880 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 881 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 882) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 883 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 884 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 885) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 886 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 887 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 888) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 889 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 890 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 891) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 892 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 893 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 894) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 895 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 896 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 897) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 898 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 899 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 900) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 901 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 902 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 903) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 904 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 905 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 906) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 907 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 908 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 909) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 910 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 911 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 912) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 913 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 914 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 915) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 916 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 917 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 918) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 919 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 920 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 921) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 922 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 923 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 924) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 925 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 926 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 927) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 928 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 929 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 930) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 931 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 932 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 933) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 934 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 935 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 936) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 937 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 938 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 939) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 940 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 941 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 942) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 943 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 944 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 945) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 946 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 947 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 948) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 949 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 950 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 951) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 952 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 953 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 954) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 955 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 956 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 957) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 958 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 959 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 960) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 961 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 962 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 963) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 964 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 965 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 966) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 967 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 968 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 969) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 970 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 971 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 972) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 973 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 974 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 975) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 976 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 977 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 978) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 979 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 980 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 981) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 982 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 983 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 984) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 985 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 986 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 987) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 988 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 989 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 990) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 991 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 992 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 993) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 994 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 995 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 996) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 997 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 998 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 999) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1000 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1001 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1002) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1003 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1004 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1005) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1006 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1007 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1008) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1009 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1010 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1011) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1012 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1013 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1014) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1015 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1016 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1017) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1018 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1019 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1020) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1021 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1022 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1023) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1024 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1025 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1026) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1027 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1028 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1029) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1030 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1031 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1032) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1033 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1034 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1035) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1036 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1037 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1038) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1039 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1040 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1041) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1042 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1043 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1044) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1045 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1046 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1047) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1048 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1049 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1050) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1051 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1052 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1053) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1054 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1055 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1056) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1057 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1058 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1059) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1060 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1061 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1062) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1063 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1064 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1065) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1066 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1067 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1068) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1069 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1070 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1071) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1072 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1073 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1074) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1075 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1076 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1077) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1078 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1079 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1080) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1081 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1082 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1083) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1084 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1085 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1086) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1087 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1088 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1089) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1090 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1091 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1092) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1093 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1094 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1095) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1096 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1097 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1098) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1099 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1100 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1101) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1102 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1103 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1104) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1105 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1106 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1107) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1108 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1109 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1110) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1111 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1112 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1113) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1114 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1115 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1116) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1117 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1118 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1119) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1120 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1121 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1122) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1123 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1124 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1125) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1126 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1127 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1128) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1129 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1130 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1131) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1132 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1133 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1134) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1135 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1136 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1137) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1138 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1139 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1140) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1141 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1142 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1143) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1144 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1145 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1146) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1147 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1148 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1149) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1150 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1151 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1152) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1153 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1154 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1155) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1156 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1157 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1158) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1159 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1160 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1161) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1162 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1163 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1164) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1165 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1166 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1167) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1168 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1169 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1170) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1171 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1172 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1173) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1174 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1175 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1176) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1177 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1178 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1179) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1180 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1181 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1182) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1183 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1184 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1185) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1186 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1187 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1188) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1189 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1190 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1191) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1192 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1193 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1194) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1195 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1196 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1197) ? o_rdata_lambda:
				    /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1198 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/
				    (r_state == zStateEstimate) &(r_counter == 1199 ) ? o_rdata_alpha:
					      /**/
					      /**/
				    /**/ 
				    (r_state == zStateEstimate) & (r_counter == 1200) ? o_rdata_lambda:
				    /**/
					      /**/
				    0;
   
   
   
   //状態遷移
   always @(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  r_state <= zStateInit;
	else if (w_trans_lambdainit)
	  r_state <= zStateLambdaInit;
	else if (w_trans_betainit)
	  r_state <= zStateBetaInit;
	else if(w_trans_row | ((r_state==zStateColumn) & (r_counter == 1602) & w_o_val_column))
	  r_state <= zStateRow;
	else if(w_trans_estimate)
	  r_state <= zStateEstimate;
	else if(w_trans_column)
	  r_state <= zStateColumn;
	else
	  r_state <= r_state;
     end // always (posedge clk or negedge xrst)
   
   //行処理の動作フラグ
   always@(posedge clk or negedge xrst)
     begin
	if (!xrst)
	  r_i_val_row <= 0;
	else if (r_i_val_row)
	  r_i_val_row <= 0;
	else if (w_trans_row)
	  r_i_val_row <= 1;
	else if (r_state == zStateRow & w_o_val_row)
	  r_i_val_row <= 1;
	else
	  r_i_val_row <= r_i_val_row;
     end // always (posedge clk or negedge xrst)
   //カウンタ
   always@(posedge clk or negedge xrst)
     begin
	if (!xrst)
	  r_counter <= 0;
	else if (r_state == zStateLambdaInit)
	  begin
	     if(r_counter == 399)
	       r_counter <= 0;
	     else
	       r_counter <= r_counter+1;
	  end
	else if (r_state == zStateBetaInit)
	  begin
	     if(r_counter == 800)
	       r_counter <= 0;
	     else
	       r_counter <= r_counter + 1;
	  end
	else if (r_state == zStateRow & w_o_val_row)
	  begin
	     if (r_counter == 2402)
	       r_counter <= 0;
	     else
	       r_counter <= r_counter + 1;
	  end
	else if (r_state ==zStateEstimate)
	  begin
	     if(r_counter == 1201)
	       r_counter<= 0;
	     else
	       r_counter <=r_counter +1;
	  end
	else if (r_state == zStateColumn & w_o_val_column)
	  begin
	     if (r_counter == 1602)
	       r_counter <=0;
	     else
	       r_counter <= r_counter + 1;
	  end
	else
	  r_counter <= r_counter;
     end // always@ (posedge clk or negedge xrst)

   //行処理の値の初期化
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  i_init_row <= 0;
	else if (i_init_row == 2 | w_trans_row==1)
	  i_init_row <=0;
	else
	  i_init_row <= i_init_row+1;
     end

   //列処理の値の初期化
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  i_init_column <= 0;
	else if ((i_init_column == 1 & r_state == zStateColumn)| w_trans_column==1 | w_trans_estimate==1 | (i_init_column == 2 & r_state== zStateEstimate))
	  i_init_column <=0;
	else
	  i_init_column <= i_init_column+1;
     end

   //繰り返し回数の更新
   always@(posedge clk or negedge xrst)
     begin
	if(!xrst)
	  r_loop <= 0;
	else if (w_trans_column)
	  r_loop <=r_loop+1;
	else
	  r_loop <= r_loop;
     end

 
   row row(
	   .i_data (o_rdata_beta[15:0]),
	   .i_val (i_val),
	   .o_data (o_data_test_alpha[15:0]),
	   .o_val (w_o_val_row),
	   .clk (clk),
	   .xrst (xrst),
	   .i_init (i_init_row [2:0])
	   );
   add add(
	   .i_data (o_column_data[15:0]),
	   .i_val (i_val),
	   .o_data (o_data_test_beta[15:0]),
	   .o_val (w_o_val_column),
	   .clk (clk),
	   .xrst (xrst),
	   .i_init (i_init_column[2:0])
	   );

   

   sram_lambda sramlambda(
	     .clk(clk),
	     .i_wen(i_wen_lambda),
	     .i_waddr(i_waddr_lambda[19:0]),
	     .i_raddr(i_raddr_lambda[19:0]),
	     .i_wdata(i_wdata_lambda[15:0]),
	     .o_rdata(o_rdata_lambda[15:0])
	     );
   sram sramalpha(
	     .clk(clk),
	     .i_wen(i_wen_alpha),
	     .i_waddr(i_waddr_alpha[19:0]),
	     .i_raddr(i_raddr_alpha[19:0]),
	     .i_wdata(i_wdata_alpha[15:0]),
	     .o_rdata(o_rdata_alpha[15:0])
	     );
   sram srambeta(
	     .clk(clk),
	     .i_wen(i_wen_beta),
	     .i_waddr(i_waddr_beta[19:0]),
	     .i_raddr(i_raddr_beta[19:0]),
	     .i_wdata(i_wdata_beta[15:0]),
	     .o_rdata(o_rdata_beta[15:0])
	     );
   
   
   
endmodule
   
	   
   
   
   

   
